
module imp_ASCON ( clk, rst, en_c, ld_rec, MuxSel1, MuxSel2, roundsel, rand_in, 
        IDt, IDst, key, DtSel, pdi_data, pdi_valid, pdi_ready, sdi_valid, 
        sdi_ready, do_data, do_ready, do_valid, rand_out );
  input [1:0] MuxSel1;
  input [63:0] rand_in;
  input [63:0] IDt;
  input [63:0] IDst;
  input [127:0] key;
  input [31:0] pdi_data;
  output [31:0] do_data;
  input [63:0] rand_out;
  input clk, rst, en_c, ld_rec, MuxSel2, roundsel, DtSel, pdi_valid, sdi_valid,
         do_ready;
  output pdi_ready, sdi_ready, do_valid;
  wire   Inst_AEAD_cmd_rd_ready, Inst_AEAD_cmd_rd_valid,
         Inst_AEAD_msg_auth_valid, Inst_AEAD_msg_auth_done,
         Inst_AEAD_bdo_ready, Inst_AEAD_bdo_valid, Inst_AEAD_cmd_wr_ready,
         Inst_AEAD_bdi_eot, Inst_AEAD_bdi_valid, Inst_AEAD_decrypt,
         Inst_AEAD_key_update, Inst_counter_n195, Inst_counter_n194,
         Inst_counter_n193, Inst_counter_n192, Inst_counter_n191,
         Inst_counter_n190, Inst_counter_n189, Inst_counter_n188,
         Inst_counter_n187, Inst_counter_n186, Inst_counter_n185,
         Inst_counter_n184, Inst_counter_n183, Inst_counter_n182,
         Inst_counter_n181, Inst_counter_n180, Inst_counter_n179,
         Inst_counter_n178, Inst_counter_n177, Inst_counter_n176,
         Inst_counter_n175, Inst_counter_n174, Inst_counter_n173,
         Inst_counter_n172, Inst_counter_n171, Inst_counter_n170,
         Inst_counter_n169, Inst_counter_n168, Inst_counter_n167,
         Inst_counter_n166, Inst_counter_n165, Inst_counter_n164,
         Inst_counter_n163, Inst_counter_n162, Inst_counter_n161,
         Inst_counter_n160, Inst_counter_n159, Inst_counter_n158,
         Inst_counter_n157, Inst_counter_n156, Inst_counter_n155,
         Inst_counter_n154, Inst_counter_n153, Inst_counter_n152,
         Inst_counter_n151, Inst_counter_n150, Inst_counter_n149,
         Inst_counter_n148, Inst_counter_n147, Inst_counter_n146,
         Inst_counter_n145, Inst_counter_n144, Inst_counter_n143,
         Inst_counter_n142, Inst_counter_n141, Inst_counter_n140,
         Inst_counter_n139, Inst_counter_n138, Inst_counter_n137,
         Inst_counter_n136, Inst_counter_n135, Inst_counter_n134,
         Inst_counter_n133, Inst_counter_n132, Inst_counter_N66,
         Inst_counter_N65, Inst_counter_N64, Inst_counter_N63,
         Inst_counter_N62, Inst_counter_N61, Inst_counter_N60,
         Inst_counter_N59, Inst_counter_N58, Inst_counter_N57,
         Inst_counter_N56, Inst_counter_N55, Inst_counter_N54,
         Inst_counter_N53, Inst_counter_N52, Inst_counter_N51,
         Inst_counter_N50, Inst_counter_N49, Inst_counter_N48,
         Inst_counter_N47, Inst_counter_N46, Inst_counter_N45,
         Inst_counter_N44, Inst_counter_N43, Inst_counter_N42,
         Inst_counter_N41, Inst_counter_N40, Inst_counter_N39,
         Inst_counter_N38, Inst_counter_N37, Inst_counter_N36,
         Inst_counter_N35, Inst_counter_N34, Inst_counter_N33,
         Inst_counter_N32, Inst_counter_N31, Inst_counter_N30,
         Inst_counter_N29, Inst_counter_N28, Inst_counter_N27,
         Inst_counter_N26, Inst_counter_N25, Inst_counter_N24,
         Inst_counter_N23, Inst_counter_N22, Inst_counter_N21,
         Inst_counter_N20, Inst_counter_N19, Inst_counter_N18,
         Inst_counter_N17, Inst_counter_N16, Inst_counter_N15,
         Inst_counter_N14, Inst_counter_N13, Inst_counter_N12,
         Inst_counter_N11, Inst_counter_N10, Inst_counter_N9, Inst_counter_N8,
         Inst_counter_N7, Inst_counter_N6, Inst_counter_N5, Inst_RegIDt_n130,
         Inst_RegIDt_n127, Inst_RegIDt_n125, Inst_RegIDt_n123,
         Inst_RegIDt_n121, Inst_RegIDt_n119, Inst_RegIDt_n117,
         Inst_RegIDt_n115, Inst_RegIDt_n113, Inst_RegIDt_n111,
         Inst_RegIDt_n109, Inst_RegIDt_n107, Inst_RegIDt_n105,
         Inst_RegIDt_n103, Inst_RegIDt_n101, Inst_RegIDt_n99, Inst_RegIDt_n97,
         Inst_RegIDt_n95, Inst_RegIDt_n93, Inst_RegIDt_n91, Inst_RegIDt_n89,
         Inst_RegIDt_n87, Inst_RegIDt_n85, Inst_RegIDt_n83, Inst_RegIDt_n81,
         Inst_RegIDt_n79, Inst_RegIDt_n77, Inst_RegIDt_n75, Inst_RegIDt_n73,
         Inst_RegIDt_n71, Inst_RegIDt_n69, Inst_RegIDt_n67, Inst_RegIDt_n65,
         Inst_RegIDt_n63, Inst_RegIDt_n61, Inst_RegIDt_n59, Inst_RegIDt_n57,
         Inst_RegIDt_n55, Inst_RegIDt_n53, Inst_RegIDt_n51, Inst_RegIDt_n49,
         Inst_RegIDt_n47, Inst_RegIDt_n45, Inst_RegIDt_n43, Inst_RegIDt_n41,
         Inst_RegIDt_n39, Inst_RegIDt_n37, Inst_RegIDt_n35, Inst_RegIDt_n33,
         Inst_RegIDt_n31, Inst_RegIDt_n29, Inst_RegIDt_n27, Inst_RegIDt_n25,
         Inst_RegIDt_n23, Inst_RegIDt_n21, Inst_RegIDt_n19, Inst_RegIDt_n17,
         Inst_RegIDt_n15, Inst_RegIDt_n13, Inst_RegIDt_n11, Inst_RegIDt_n9,
         Inst_RegIDt_n7, Inst_RegIDt_n5, Inst_RegIDt_n3,
         Inst_AEAD_u_input_n554, Inst_AEAD_u_input_n553,
         Inst_AEAD_u_input_n552, Inst_AEAD_u_input_n551,
         Inst_AEAD_u_input_n550, Inst_AEAD_u_input_n549,
         Inst_AEAD_u_input_n548, Inst_AEAD_u_input_n547,
         Inst_AEAD_u_input_n546, Inst_AEAD_u_input_n545,
         Inst_AEAD_u_input_n544, Inst_AEAD_u_input_n543,
         Inst_AEAD_u_input_n542, Inst_AEAD_u_input_n541,
         Inst_AEAD_u_input_n540, Inst_AEAD_u_input_n539,
         Inst_AEAD_u_input_n538, Inst_AEAD_u_input_n537,
         Inst_AEAD_u_input_n536, Inst_AEAD_u_input_n535,
         Inst_AEAD_u_input_n534, Inst_AEAD_u_input_n533,
         Inst_AEAD_u_input_n532, Inst_AEAD_u_input_n531,
         Inst_AEAD_u_input_n530, Inst_AEAD_u_input_n529,
         Inst_AEAD_u_input_n528, Inst_AEAD_u_input_n527,
         Inst_AEAD_u_input_n526, Inst_AEAD_u_input_n525,
         Inst_AEAD_u_input_n524, Inst_AEAD_u_input_n523,
         Inst_AEAD_u_input_n522, Inst_AEAD_u_input_n521,
         Inst_AEAD_u_input_n520, Inst_AEAD_u_input_n519,
         Inst_AEAD_u_input_n518, Inst_AEAD_u_input_n517,
         Inst_AEAD_u_input_n516, Inst_AEAD_u_input_n515,
         Inst_AEAD_u_input_n514, Inst_AEAD_u_input_n513,
         Inst_AEAD_u_input_n512, Inst_AEAD_u_input_n511,
         Inst_AEAD_u_input_n510, Inst_AEAD_u_input_n509,
         Inst_AEAD_u_input_n508, Inst_AEAD_u_input_n507,
         Inst_AEAD_u_input_n506, Inst_AEAD_u_input_n505,
         Inst_AEAD_u_input_n504, Inst_AEAD_u_input_n503,
         Inst_AEAD_u_input_n502, Inst_AEAD_u_input_n501,
         Inst_AEAD_u_input_n500, Inst_AEAD_u_input_n499,
         Inst_AEAD_u_input_n498, Inst_AEAD_u_input_n497,
         Inst_AEAD_u_input_n496, Inst_AEAD_u_input_n495,
         Inst_AEAD_u_input_n494, Inst_AEAD_u_input_n493,
         Inst_AEAD_u_input_n492, Inst_AEAD_u_input_n491,
         Inst_AEAD_u_input_n490, Inst_AEAD_u_input_n489,
         Inst_AEAD_u_input_n488, Inst_AEAD_u_input_n487,
         Inst_AEAD_u_input_n486, Inst_AEAD_u_input_n485,
         Inst_AEAD_u_input_n484, Inst_AEAD_u_input_n483,
         Inst_AEAD_u_input_n482, Inst_AEAD_u_input_n481,
         Inst_AEAD_u_input_n480, Inst_AEAD_u_input_n479,
         Inst_AEAD_u_input_n478, Inst_AEAD_u_input_n477,
         Inst_AEAD_u_input_n421, Inst_AEAD_u_input_n392,
         Inst_AEAD_u_input_n391, Inst_AEAD_u_input_n362,
         Inst_AEAD_u_input_n358, Inst_AEAD_u_input_n321,
         Inst_AEAD_u_input_n320, Inst_AEAD_u_input_n319,
         Inst_AEAD_u_input_n318, Inst_AEAD_u_input_n317,
         Inst_AEAD_u_input_n316, Inst_AEAD_u_input_n315,
         Inst_AEAD_u_input_n314, Inst_AEAD_u_input_n313,
         Inst_AEAD_u_input_n312, Inst_AEAD_u_input_n311,
         Inst_AEAD_u_input_n310, Inst_AEAD_u_input_n309,
         Inst_AEAD_u_input_n308, Inst_AEAD_u_input_n307,
         Inst_AEAD_u_input_n306, Inst_AEAD_u_input_n305,
         Inst_AEAD_u_input_n304, Inst_AEAD_u_input_n303,
         Inst_AEAD_u_input_n287, Inst_AEAD_u_input_n286, Inst_AEAD_u_input_n85,
         Inst_AEAD_u_input_ctr_0_, Inst_AEAD_u_input_is_extra,
         Inst_AEAD_u_input_N220, Inst_AEAD_u_input_N219,
         Inst_AEAD_u_input_N218, Inst_AEAD_u_input_N217,
         Inst_AEAD_u_input_slen_1_, Inst_AEAD_u_input_slen_2_,
         Inst_AEAD_u_input_slen_3_, Inst_AEAD_u_input_slen_4_,
         Inst_AEAD_u_input_slen_5_, Inst_AEAD_u_input_slen_6_,
         Inst_AEAD_u_input_N143, Inst_AEAD_u_input_N142,
         Inst_AEAD_u_input_N141, Inst_AEAD_u_input_N140,
         Inst_AEAD_u_input_N139, Inst_AEAD_u_input_N138,
         Inst_AEAD_u_input_N137, Inst_AEAD_u_input_N136,
         Inst_AEAD_u_input_N135, Inst_AEAD_u_input_N134,
         Inst_AEAD_u_input_N133, Inst_AEAD_u_input_N132,
         Inst_AEAD_u_input_N131, Inst_AEAD_u_input_N128,
         Inst_AEAD_u_input_sgmt_len_1_, Inst_AEAD_u_input_sgmt_len_2_,
         Inst_AEAD_u_input_sgmt_len_3_, Inst_AEAD_u_input_sgmt_len_4_,
         Inst_AEAD_u_input_sgmt_len_5_, Inst_AEAD_u_input_sgmt_len_6_,
         Inst_AEAD_u_input_sgmt_len_7_, Inst_AEAD_u_input_sgmt_len_8_,
         Inst_AEAD_u_input_sgmt_len_9_, Inst_AEAD_u_input_sgmt_len_10_,
         Inst_AEAD_u_input_sgmt_len_11_, Inst_AEAD_u_input_sgmt_len_12_,
         Inst_AEAD_u_input_sgmt_len_13_, Inst_AEAD_u_input_sgmt_len_14_,
         Inst_AEAD_u_input_sgmt_len_15_, Inst_AEAD_u_input_ss_0_,
         Inst_AEAD_u_input_ss_1_, Inst_AEAD_u_input_ps_0_,
         Inst_AEAD_u_input_ps_1_, Inst_AEAD_u_input_ps_2_,
         Inst_AEAD_u_input_size_0_, Inst_AEAD_u_input_size_1_,
         Inst_AEAD_u_input_vbytes_3_, Inst_AEAD_u_input_req_pad,
         Inst_AEAD_u_input_ploc_0_, Inst_AEAD_u_input_ploc_1_,
         Inst_AEAD_u_input_reg_sel_zero, Inst_AEAD_u_cc_sel_key_lo,
         Inst_AEAD_u_cc_en_cmp, Inst_AEAD_u_cc_en_state,
         Inst_AEAD_u_hdr_buffer_n435, Inst_AEAD_u_hdr_buffer_n434,
         Inst_AEAD_u_hdr_buffer_n433, Inst_AEAD_u_hdr_buffer_n432,
         Inst_AEAD_u_hdr_buffer_n431, Inst_AEAD_u_hdr_buffer_n430,
         Inst_AEAD_u_hdr_buffer_n429, Inst_AEAD_u_hdr_buffer_n428,
         Inst_AEAD_u_hdr_buffer_n427, Inst_AEAD_u_hdr_buffer_n426,
         Inst_AEAD_u_hdr_buffer_n424, Inst_AEAD_u_hdr_buffer_n423,
         Inst_AEAD_u_hdr_buffer_n422, Inst_AEAD_u_hdr_buffer_n421,
         Inst_AEAD_u_hdr_buffer_n420, Inst_AEAD_u_hdr_buffer_n419,
         Inst_AEAD_u_hdr_buffer_n418, Inst_AEAD_u_hdr_buffer_n417,
         Inst_AEAD_u_hdr_buffer_n416, Inst_AEAD_u_hdr_buffer_n415,
         Inst_AEAD_u_hdr_buffer_n414, Inst_AEAD_u_hdr_buffer_n413,
         Inst_AEAD_u_hdr_buffer_n412, Inst_AEAD_u_hdr_buffer_n411,
         Inst_AEAD_u_hdr_buffer_n410, Inst_AEAD_u_hdr_buffer_n409,
         Inst_AEAD_u_hdr_buffer_n408, Inst_AEAD_u_hdr_buffer_n407,
         Inst_AEAD_u_hdr_buffer_n406, Inst_AEAD_u_hdr_buffer_n405,
         Inst_AEAD_u_hdr_buffer_n404, Inst_AEAD_u_hdr_buffer_n403,
         Inst_AEAD_u_hdr_buffer_n402, Inst_AEAD_u_hdr_buffer_n400,
         Inst_AEAD_u_hdr_buffer_n399, Inst_AEAD_u_hdr_buffer_n398,
         Inst_AEAD_u_hdr_buffer_n397, Inst_AEAD_u_hdr_buffer_n396,
         Inst_AEAD_u_hdr_buffer_n395, Inst_AEAD_u_hdr_buffer_n394,
         Inst_AEAD_u_hdr_buffer_n393, Inst_AEAD_u_hdr_buffer_n392,
         Inst_AEAD_u_hdr_buffer_n391, Inst_AEAD_u_hdr_buffer_n390,
         Inst_AEAD_u_hdr_buffer_n389, Inst_AEAD_u_hdr_buffer_n388,
         Inst_AEAD_u_hdr_buffer_n387, Inst_AEAD_u_hdr_buffer_n386,
         Inst_AEAD_u_hdr_buffer_n385, Inst_AEAD_u_hdr_buffer_n384,
         Inst_AEAD_u_hdr_buffer_n383, Inst_AEAD_u_hdr_buffer_n374,
         Inst_AEAD_u_hdr_buffer_n326, Inst_AEAD_u_hdr_buffer_n294,
         Inst_AEAD_u_hdr_buffer_n293, Inst_AEAD_u_hdr_buffer_n292,
         Inst_AEAD_u_hdr_buffer_n291, Inst_AEAD_u_hdr_buffer_n290,
         Inst_AEAD_u_hdr_buffer_n289, Inst_AEAD_u_hdr_buffer_n288,
         Inst_AEAD_u_hdr_buffer_n287, Inst_AEAD_u_hdr_buffer_n286,
         Inst_AEAD_u_hdr_buffer_n285, Inst_AEAD_u_hdr_buffer_n284,
         Inst_AEAD_u_hdr_buffer_n283, Inst_AEAD_u_hdr_buffer_n282,
         Inst_AEAD_u_hdr_buffer_n281, Inst_AEAD_u_hdr_buffer_n280,
         Inst_AEAD_u_hdr_buffer_n279, Inst_AEAD_u_hdr_buffer_n278,
         Inst_AEAD_u_hdr_buffer_n277, Inst_AEAD_u_hdr_buffer_n276,
         Inst_AEAD_u_hdr_buffer_n275, Inst_AEAD_u_hdr_buffer_n274,
         Inst_AEAD_u_hdr_buffer_n273, Inst_AEAD_u_hdr_buffer_n272,
         Inst_AEAD_u_hdr_buffer_n271, Inst_AEAD_u_hdr_buffer_N366,
         Inst_AEAD_u_hdr_buffer_N365, Inst_AEAD_u_hdr_buffer_N364,
         Inst_AEAD_u_hdr_buffer_N363, Inst_AEAD_u_hdr_buffer_N362,
         Inst_AEAD_u_hdr_buffer_N361, Inst_AEAD_u_hdr_buffer_N360,
         Inst_AEAD_u_hdr_buffer_N359, Inst_AEAD_u_hdr_buffer_N358,
         Inst_AEAD_u_hdr_buffer_N357, Inst_AEAD_u_hdr_buffer_N356,
         Inst_AEAD_u_hdr_buffer_N355, Inst_AEAD_u_hdr_buffer_N354,
         Inst_AEAD_u_hdr_buffer_N353, Inst_AEAD_u_hdr_buffer_N352,
         Inst_AEAD_u_hdr_buffer_N351, Inst_AEAD_u_hdr_buffer_N350,
         Inst_AEAD_u_hdr_buffer_N349, Inst_AEAD_u_hdr_buffer_N348,
         Inst_AEAD_u_hdr_buffer_N347, Inst_AEAD_u_hdr_buffer_N346,
         Inst_AEAD_u_hdr_buffer_N345, Inst_AEAD_u_hdr_buffer_N344,
         Inst_AEAD_u_hdr_buffer_N343, Inst_AEAD_u_hdr_buffer_memory_0__0_,
         Inst_AEAD_u_hdr_buffer_memory_0__1_,
         Inst_AEAD_u_hdr_buffer_memory_0__2_,
         Inst_AEAD_u_hdr_buffer_memory_0__3_,
         Inst_AEAD_u_hdr_buffer_memory_0__4_,
         Inst_AEAD_u_hdr_buffer_memory_0__5_,
         Inst_AEAD_u_hdr_buffer_memory_0__6_,
         Inst_AEAD_u_hdr_buffer_memory_0__7_,
         Inst_AEAD_u_hdr_buffer_memory_0__8_,
         Inst_AEAD_u_hdr_buffer_memory_0__9_,
         Inst_AEAD_u_hdr_buffer_memory_0__10_,
         Inst_AEAD_u_hdr_buffer_memory_0__11_,
         Inst_AEAD_u_hdr_buffer_memory_0__12_,
         Inst_AEAD_u_hdr_buffer_memory_0__13_,
         Inst_AEAD_u_hdr_buffer_memory_0__14_,
         Inst_AEAD_u_hdr_buffer_memory_0__15_,
         Inst_AEAD_u_hdr_buffer_memory_0__16_,
         Inst_AEAD_u_hdr_buffer_memory_0__17_,
         Inst_AEAD_u_hdr_buffer_memory_0__18_,
         Inst_AEAD_u_hdr_buffer_memory_0__19_,
         Inst_AEAD_u_hdr_buffer_memory_0__20_,
         Inst_AEAD_u_hdr_buffer_memory_0__21_,
         Inst_AEAD_u_hdr_buffer_memory_0__22_,
         Inst_AEAD_u_hdr_buffer_memory_0__23_,
         Inst_AEAD_u_hdr_buffer_memory_1__0_,
         Inst_AEAD_u_hdr_buffer_memory_1__1_,
         Inst_AEAD_u_hdr_buffer_memory_1__2_,
         Inst_AEAD_u_hdr_buffer_memory_1__3_,
         Inst_AEAD_u_hdr_buffer_memory_1__4_,
         Inst_AEAD_u_hdr_buffer_memory_1__5_,
         Inst_AEAD_u_hdr_buffer_memory_1__6_,
         Inst_AEAD_u_hdr_buffer_memory_1__7_,
         Inst_AEAD_u_hdr_buffer_memory_1__8_,
         Inst_AEAD_u_hdr_buffer_memory_1__9_,
         Inst_AEAD_u_hdr_buffer_memory_1__10_,
         Inst_AEAD_u_hdr_buffer_memory_1__11_,
         Inst_AEAD_u_hdr_buffer_memory_1__12_,
         Inst_AEAD_u_hdr_buffer_memory_1__13_,
         Inst_AEAD_u_hdr_buffer_memory_1__14_,
         Inst_AEAD_u_hdr_buffer_memory_1__15_,
         Inst_AEAD_u_hdr_buffer_memory_1__16_,
         Inst_AEAD_u_hdr_buffer_memory_1__17_,
         Inst_AEAD_u_hdr_buffer_memory_1__18_,
         Inst_AEAD_u_hdr_buffer_memory_1__19_,
         Inst_AEAD_u_hdr_buffer_memory_1__20_,
         Inst_AEAD_u_hdr_buffer_memory_1__21_,
         Inst_AEAD_u_hdr_buffer_memory_1__22_,
         Inst_AEAD_u_hdr_buffer_memory_1__23_,
         Inst_AEAD_u_hdr_buffer_memory_2__0_,
         Inst_AEAD_u_hdr_buffer_memory_2__1_,
         Inst_AEAD_u_hdr_buffer_memory_2__2_,
         Inst_AEAD_u_hdr_buffer_memory_2__3_,
         Inst_AEAD_u_hdr_buffer_memory_2__4_,
         Inst_AEAD_u_hdr_buffer_memory_2__5_,
         Inst_AEAD_u_hdr_buffer_memory_2__6_,
         Inst_AEAD_u_hdr_buffer_memory_2__7_,
         Inst_AEAD_u_hdr_buffer_memory_2__8_,
         Inst_AEAD_u_hdr_buffer_memory_2__9_,
         Inst_AEAD_u_hdr_buffer_memory_2__10_,
         Inst_AEAD_u_hdr_buffer_memory_2__11_,
         Inst_AEAD_u_hdr_buffer_memory_2__12_,
         Inst_AEAD_u_hdr_buffer_memory_2__13_,
         Inst_AEAD_u_hdr_buffer_memory_2__14_,
         Inst_AEAD_u_hdr_buffer_memory_2__15_,
         Inst_AEAD_u_hdr_buffer_memory_2__16_,
         Inst_AEAD_u_hdr_buffer_memory_2__17_,
         Inst_AEAD_u_hdr_buffer_memory_2__18_,
         Inst_AEAD_u_hdr_buffer_memory_2__19_,
         Inst_AEAD_u_hdr_buffer_memory_2__20_,
         Inst_AEAD_u_hdr_buffer_memory_2__21_,
         Inst_AEAD_u_hdr_buffer_memory_2__22_,
         Inst_AEAD_u_hdr_buffer_memory_2__23_, Inst_AEAD_u_hdr_buffer_looped,
         Inst_AEAD_u_hdr_buffer_wrptr_0_, Inst_AEAD_u_hdr_buffer_wrptr_1_,
         Inst_AEAD_u_cc_u_cc_dp_n2204, Inst_AEAD_u_cc_u_cc_dp_n2203,
         Inst_AEAD_u_cc_u_cc_dp_n2202, Inst_AEAD_u_cc_u_cc_dp_n2201,
         Inst_AEAD_u_cc_u_cc_dp_n2200, Inst_AEAD_u_cc_u_cc_dp_n2199,
         Inst_AEAD_u_cc_u_cc_dp_N712, Inst_AEAD_u_cc_u_cc_dp_rc_0_,
         Inst_AEAD_u_cc_u_cc_dp_rc_1_, Inst_AEAD_u_cc_u_cc_dp_rc_2_,
         Inst_AEAD_u_cc_u_cc_dp_rc_3_, Inst_AEAD_u_cc_u_cc_dp_rc_4_,
         Inst_AEAD_u_cc_u_cc_dp_rc_5_, Inst_AEAD_u_cc_u_cc_dp_rc_6_,
         Inst_AEAD_u_cc_u_cc_dp_rc_7_, Inst_AEAD_u_cc_u_cc_dp_reg_key_0_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_1_, Inst_AEAD_u_cc_u_cc_dp_reg_key_2_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_3_, Inst_AEAD_u_cc_u_cc_dp_reg_key_4_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_5_, Inst_AEAD_u_cc_u_cc_dp_reg_key_6_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_7_, Inst_AEAD_u_cc_u_cc_dp_reg_key_8_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_9_, Inst_AEAD_u_cc_u_cc_dp_reg_key_10_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_11_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_12_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_13_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_14_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_15_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_16_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_17_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_18_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_19_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_20_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_21_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_22_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_23_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_24_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_25_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_26_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_27_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_28_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_29_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_30_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_31_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_32_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_33_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_34_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_35_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_36_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_37_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_38_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_39_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_40_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_41_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_42_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_43_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_44_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_45_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_46_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_47_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_48_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_49_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_50_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_51_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_52_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_53_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_54_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_55_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_56_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_57_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_58_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_59_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_60_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_61_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_62_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_63_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_64_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_65_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_66_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_67_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_68_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_69_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_70_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_71_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_72_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_73_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_74_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_75_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_76_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_77_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_78_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_79_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_80_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_81_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_82_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_83_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_84_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_85_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_86_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_87_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_88_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_89_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_90_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_91_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_92_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_93_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_94_,
         Inst_AEAD_u_cc_u_cc_dp_reg_key_95_, Inst_AEAD_u_cc_u_cc_ctrl_n123,
         Inst_AEAD_u_cc_u_cc_ctrl_n122, Inst_AEAD_u_cc_u_cc_ctrl_n121,
         Inst_AEAD_u_cc_u_cc_ctrl_n120, Inst_AEAD_u_cc_u_cc_ctrl_n119,
         Inst_AEAD_u_cc_u_cc_ctrl_n118, Inst_AEAD_u_cc_u_cc_ctrl_n117,
         Inst_AEAD_u_cc_u_cc_ctrl_n116, Inst_AEAD_u_cc_u_cc_ctrl_n115,
         Inst_AEAD_u_cc_u_cc_ctrl_n114, Inst_AEAD_u_cc_u_cc_ctrl_n113,
         Inst_AEAD_u_cc_u_cc_ctrl_n112, Inst_AEAD_u_cc_u_cc_ctrl_n52,
         Inst_AEAD_u_cc_u_cc_ctrl_n37, Inst_AEAD_u_cc_u_cc_ctrl_is_init_dat,
         Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_1_,
         Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_2_,
         Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_3_, Inst_AEAD_u_cc_u_cc_ctrl_state_0_,
         Inst_AEAD_u_cc_u_cc_ctrl_state_1_, Inst_AEAD_u_cc_u_cc_ctrl_state_2_,
         Inst_AEAD_u_cc_u_cc_ctrl_round_1_, Inst_AEAD_u_cc_u_cc_ctrl_round_2_,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5088, n5090, n5092, n5094, n5096, n5098,
         n5100, n5102, n5104, n5106, n5108, n5110, n5112, n5114, n5116, n5118,
         n5120, n5122, n5124, n5126, n5128, n5130, n5132, n5134, n5136, n5138,
         n5140, n5142, n5144, n5146, n5148, n5150, n5152, n5154, n5156, n5158,
         n5160, n5162, n5164, n5166, n5168, n5170, n5172, n5174, n5176, n5178,
         n5180, n5182, n5184, n5186, n5188, n5190, n5192, n5194, n5196, n5198,
         n5200, n5202, n5204, n5206, n5208, n5210, n5212, n5214;
  wire   [63:0] randd;
  wire   [63:0] IDtReg;
  wire   [63:0] IDstReg;
  wire   [23:0] Inst_AEAD_cmd_dout;
  wire   [63:0] Inst_AEAD_bdo;
  wire   [7:0] Inst_AEAD_bdi_valid_bytes;
  wire   [3:0] Inst_AEAD_bdi_size;
  wire   [63:0] Inst_AEAD_bdi;
  wire   [31:0] Inst_AEAD_key;
  wire   [1:0] Inst_AEAD_u_cc_sel_tag;
  wire   [319:0] Inst_AEAD_u_cc_u_cc_dp_istate;
  wire   [15:4] Inst_AEAD_u_input_sub_751_carry;
  wire   [6:4] Inst_AEAD_u_input_sub_774_carry;
  wire   [63:2] Inst_counter_add_3021_carry;

  PostProcessor Inst_AEAD_u_output ( .clk(clk), .rst(rst), .do_data(do_data), 
        .do_ready(do_ready), .do_valid(do_valid), .cmd(Inst_AEAD_cmd_dout), 
        .cmd_valid(Inst_AEAD_cmd_rd_valid), .cmd_ready(Inst_AEAD_cmd_rd_ready), 
        .bdo(Inst_AEAD_bdo), .bdo_valid(Inst_AEAD_bdo_valid), .bdo_ready(
        Inst_AEAD_bdo_ready), .bdo_size({1'b0, 1'b0, 1'b0, 1'b0}), 
        .msg_auth_done(Inst_AEAD_msg_auth_done), .msg_auth_valid(
        Inst_AEAD_msg_auth_valid) );
  SEDFFXL Inst_AEAD_u_input_size_reg_2_ ( .D(n5085), .SI(1'b0), .E(
        Inst_AEAD_u_input_n392), .SE(1'b0), .CK(clk), .QN(n1567) );
  SEDFFXL Inst_AEAD_u_input_sgmt_lst_reg ( .D(pdi_data[24]), .SI(1'b0), .E(
        Inst_AEAD_u_input_n554), .SE(1'b0), .CK(clk), .QN(n1566) );
  SEDFFXL Inst_AEAD_u_input_sgmt_type_reg_3_ ( .D(pdi_data[31]), .SI(1'b0), 
        .E(Inst_AEAD_u_input_n554), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_input_n358) );
  SEDFFXL Inst_AEAD_u_input_sgmt_type_reg_2_ ( .D(pdi_data[30]), .SI(1'b0), 
        .E(Inst_AEAD_u_input_n554), .SE(1'b0), .CK(clk), .Q(n468), .QN(n1564)
         );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__0_ ( .D(pdi_data[0]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n294) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__1_ ( .D(pdi_data[1]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n293) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__2_ ( .D(pdi_data[2]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n292) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__3_ ( .D(pdi_data[3]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n291) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__4_ ( .D(pdi_data[4]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n290) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__5_ ( .D(pdi_data[5]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n289) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__6_ ( .D(pdi_data[6]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n288) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__7_ ( .D(pdi_data[7]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n287) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__8_ ( .D(pdi_data[8]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n286) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__9_ ( .D(pdi_data[9]), .SI(1'b0), 
        .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n285) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__10_ ( .D(pdi_data[10]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n284) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__11_ ( .D(pdi_data[11]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n283) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__12_ ( .D(pdi_data[12]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n282) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__13_ ( .D(pdi_data[13]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n281) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__14_ ( .D(pdi_data[14]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n280) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__15_ ( .D(pdi_data[15]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n279) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__16_ ( .D(pdi_data[24]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n278) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__17_ ( .D(pdi_data[25]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n277) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__18_ ( .D(1'b0), .SI(1'b0), .E(
        Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n276) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__19_ ( .D(pdi_data[27]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n275) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__20_ ( .D(pdi_data[28]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n274) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__21_ ( .D(pdi_data[29]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n273) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__22_ ( .D(pdi_data[30]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n272) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_3__23_ ( .D(pdi_data[31]), .SI(
        1'b0), .E(Inst_AEAD_u_hdr_buffer_n326), .SE(1'b0), .CK(clk), .QN(
        Inst_AEAD_u_hdr_buffer_n271) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_msg_auth_valid_r_reg ( .D(
        Inst_AEAD_u_cc_u_cc_dp_N712), .SI(1'b0), .E(Inst_AEAD_u_cc_en_cmp), 
        .SE(1'b0), .CK(clk), .QN(n1561) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_319_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[319]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1560) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_318_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[318]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n354), .QN(n1559) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_317_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[317]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .Q(n356), .QN(n1558) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_316_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[316]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .Q(n358), .QN(n1557) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_315_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[315]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .Q(n360), .QN(n1556) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_314_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[314]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .Q(n362), .QN(n1555) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_313_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[313]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .Q(n344), .QN(n1554) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_312_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[312]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n345), .QN(n1553) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_311_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[311]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n346), .QN(n1552) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_310_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[310]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1551) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_309_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[309]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .Q(n347), .QN(n1550) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_308_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[308]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n359), .QN(n1549) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_307_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[307]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n361), .QN(n1548) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_306_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[306]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .Q(n364), .QN(n1547) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_305_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[305]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .Q(n365), .QN(n1546) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_304_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[304]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .Q(n366), .QN(n1545) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_303_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[303]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .Q(n367), .QN(n1544) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_302_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[302]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .Q(n369), .QN(n1543) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_301_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[301]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .Q(n355), .QN(n1542) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_300_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[300]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n357), .QN(n1541) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_299_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[299]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .Q(n379), .QN(n1540) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_298_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[298]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n380), .QN(n1539) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_297_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[297]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .Q(n370), .QN(n1538) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_296_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[296]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .Q(n363), .QN(n1537) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_295_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[295]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n351), .QN(n1536) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_294_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[294]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .Q(n352), .QN(n1535) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_293_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[293]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .Q(n353), .QN(n1534) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_292_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[292]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .Q(n368), .QN(n1533) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_291_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[291]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .Q(n374), .QN(n1532) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_290_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[290]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n342), .QN(n1531) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_289_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[289]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n343), .QN(n1530) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_288_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[288]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n375), .QN(n1529) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_287_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[287]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1528) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_286_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[286]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1527) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_285_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[285]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .QN(n1526) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_284_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[284]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .QN(n1525) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_283_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[283]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1524) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_282_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[282]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1523) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_281_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[281]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .QN(n1522) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_280_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[280]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1521) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_279_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[279]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1520) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_278_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[278]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .QN(n1519) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_277_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[277]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1518) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_276_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[276]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1517) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_275_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[275]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1516) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_274_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[274]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1515) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_273_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[273]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .QN(n1514) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_272_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[272]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n348), .QN(n1513) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_271_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[271]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .Q(n349), .QN(n1512) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_270_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[270]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n371), .QN(n1511) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_269_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[269]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1510) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_268_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[268]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1509) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_267_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[267]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1508) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_266_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[266]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1507) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_265_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[265]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .Q(n372), .QN(n1506) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_264_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[264]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n373), .QN(n1505) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_263_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[263]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n350), .QN(n1504) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_262_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[262]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .QN(n1503) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_261_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[261]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1502) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_260_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[260]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1501) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_259_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[259]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1500) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_258_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[258]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1499) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_257_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[257]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1498) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_256_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[256]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1497) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_255_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[255]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1496) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_254_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[254]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1495) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_253_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[253]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .QN(n1494) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_252_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[252]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1493) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_251_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[251]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1492) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_250_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[250]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1491) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_249_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[249]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1490) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_248_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[248]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1489) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_247_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[247]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .QN(n1488) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_246_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[246]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1487) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_245_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[245]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1486) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_244_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[244]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1485) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_243_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[243]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .QN(n1484) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_242_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[242]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1483) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_241_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[241]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1482) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_240_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[240]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1481) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_239_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[239]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1480) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_238_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[238]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1479) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_237_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[237]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .QN(n1478) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_236_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[236]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .QN(n1477) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_235_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[235]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1476) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_234_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[234]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .QN(n1475) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_233_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[233]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1474) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_232_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[232]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1473) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_231_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[231]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1472) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_230_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[230]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1471) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_229_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[229]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1470) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_228_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[228]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1469) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_227_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[227]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1468) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_226_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[226]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1467) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_225_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[225]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1466) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_224_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[224]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1465) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_223_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[223]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1464) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_222_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[222]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1463) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_221_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[221]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .QN(n1462) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_220_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[220]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .QN(n1461) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_219_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[219]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1460) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_218_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[218]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1459) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_217_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[217]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1458) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_216_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[216]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .QN(n1457) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_215_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[215]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1456) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_214_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[214]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .QN(n1455) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_213_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[213]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1454) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_212_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[212]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1453) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_211_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[211]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1452) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_210_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[210]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1451) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_209_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[209]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1450) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_208_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[208]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1449) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_207_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[207]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1448) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_206_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[206]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1447) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_205_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[205]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1446) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_204_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[204]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1445) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_203_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[203]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1444) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_202_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[202]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1443) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_201_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[201]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .QN(n1442) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_200_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[200]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1441) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_199_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[199]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n341), .QN(n1440) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_198_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[198]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1439) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_197_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[197]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1438) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_196_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[196]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1437) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_195_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[195]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1436) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_194_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[194]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1435) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_193_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[193]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1434) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_192_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[192]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1433) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_191_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[191]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1432) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_190_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[190]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1431) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_189_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[189]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1430) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_188_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[188]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1429) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_187_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[187]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1428) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_186_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[186]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1427) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_185_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[185]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1426) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_184_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[184]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1425) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_183_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[183]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1424) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_182_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[182]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1423) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_181_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[181]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1422) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_180_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[180]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1421) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_179_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[179]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .QN(n1420) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_178_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[178]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1419) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_177_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[177]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1418) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_176_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[176]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1417) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_175_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[175]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1416) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_174_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[174]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1415) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_173_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[173]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1414) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_172_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[172]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1413) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_171_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[171]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1412) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_170_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[170]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1411) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_169_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[169]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1410) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_168_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[168]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1409) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_167_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[167]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1408) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_166_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[166]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1407) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_165_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[165]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1406) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_164_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[164]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1405) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_163_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[163]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1404) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_162_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[162]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1403) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_161_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[161]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1402) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_160_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[160]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1401) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_159_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[159]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1400) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_158_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[158]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1399) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_157_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[157]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1398) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_156_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[156]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1397) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_155_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[155]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1396) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_154_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[154]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1395) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_153_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[153]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1394) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_152_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[152]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .QN(n1393) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_151_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[151]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1392) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_150_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[150]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1391) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_149_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[149]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1390) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_148_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[148]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .QN(n1389) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_147_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[147]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1388) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_146_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[146]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1387) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_145_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[145]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .QN(n1386) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_144_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[144]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1385) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_143_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[143]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .QN(n1384) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_142_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[142]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1383) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_141_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[141]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1382) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_140_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[140]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1381) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_139_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[139]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1380) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_138_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[138]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .QN(n1379) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_137_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[137]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1378) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_136_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[136]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1377) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_135_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[135]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1376) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_134_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[134]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1375) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_133_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[133]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1374) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_132_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[132]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1373) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_131_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[131]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1372) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_130_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[130]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1371) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_129_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[129]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1370) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_128_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[128]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1369) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_127_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[127]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1368) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_126_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[126]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1367) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_125_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[125]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1366) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_124_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[124]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .QN(n1365) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_123_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[123]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .QN(n1364) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_122_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[122]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .QN(n1363) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_121_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[121]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .QN(n1362) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_120_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[120]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1361) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_119_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[119]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1360) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_118_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[118]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1359) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_117_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[117]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1358) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_116_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[116]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1357) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_115_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[115]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1356) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_114_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[114]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1355) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_113_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[113]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1354) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_112_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[112]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1353) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_111_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[111]), .SI(1'b0), .E(n1018), .SE(1'b0), 
        .CK(clk), .QN(n1352) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_110_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[110]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1351) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_109_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[109]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1350) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_108_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[108]), .SI(1'b0), .E(n1002), .SE(1'b0), 
        .CK(clk), .QN(n1349) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_107_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[107]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .QN(n1348) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_106_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[106]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .QN(n1347) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_105_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[105]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .QN(n1346) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_104_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[104]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1345) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_103_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[103]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .QN(n1344) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_102_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[102]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1343) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_101_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[101]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1342) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_100_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[100]), .SI(1'b0), .E(n1009), .SE(1'b0), 
        .CK(clk), .QN(n1341) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_99_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[99]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .Q(n445), .QN(n1340) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_98_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[98]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n446), .QN(n1339) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_97_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[97]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n447), .QN(n1338) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_96_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[96]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n448), .QN(n1337) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_95_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[95]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .Q(n449), .QN(n1336) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_94_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[94]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .Q(n450), .QN(n1335) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_93_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[93]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n451), .QN(n1334) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_92_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[92]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .Q(n452), .QN(n1333) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_91_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[91]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .Q(n453), .QN(n1332) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_90_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[90]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .Q(n454), .QN(n1331) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_89_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[89]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n455), .QN(n1330) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_88_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[88]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .Q(n456), .QN(n1329) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_87_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[87]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .Q(n457), .QN(n1328) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_86_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[86]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .Q(n458), .QN(n1327) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_85_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[85]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .Q(n459), .QN(n1326) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_84_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[84]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n443), .QN(n1325) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_83_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[83]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .Q(n444), .QN(n1324) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_82_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[82]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .Q(n463), .QN(n1323) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_81_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[81]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n465), .QN(n1322) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_80_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[80]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1321) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_79_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[79]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .QN(n1320) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_78_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[78]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .QN(n1319) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_77_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[77]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .Q(n460), .QN(n1318) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_76_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[76]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n461), .QN(n1317) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_75_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[75]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .Q(n462), .QN(n1316) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_74_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[74]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n464), .QN(n1315) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_73_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[73]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .QN(n1314) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_72_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[72]), .SI(1'b0), .E(n1019), .SE(1'b0), 
        .CK(clk), .QN(n1313) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_71_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[71]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n441), .QN(n1312) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_70_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[70]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .Q(n435), .QN(n1311) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_69_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[69]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n436), .QN(n1310) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_68_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[68]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .Q(n437), .QN(n1309) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_67_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[67]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .Q(n438), .QN(n1308) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_66_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[66]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .Q(n439), .QN(n1307) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_65_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[65]), .SI(1'b0), .E(n1003), .SE(1'b0), 
        .CK(clk), .Q(n440), .QN(n1306) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_63_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[63]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .Q(n381), .QN(n1305) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_62_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[62]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n382), .QN(n1304) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_61_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[61]), .SI(1'b0), .E(n1028), .SE(1'b0), 
        .CK(clk), .Q(n383), .QN(n1303) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_60_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[60]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .Q(n384), .QN(n1302) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_59_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[59]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .Q(n385), .QN(n1301) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_58_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[58]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .Q(n386), .QN(n1300) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_57_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[57]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .Q(n387), .QN(n1299) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_56_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[56]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .Q(n388), .QN(n1298) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_55_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[55]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .Q(n389), .QN(n1297) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_54_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[54]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .Q(n390), .QN(n1296) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_53_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[53]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .Q(n391), .QN(n1295) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_52_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[52]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n392), .QN(n1294) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_51_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[51]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n393), .QN(n1293) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_50_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[50]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .Q(n394), .QN(n1292) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_49_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[49]), .SI(1'b0), .E(n1022), .SE(1'b0), 
        .CK(clk), .Q(n395), .QN(n1291) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_48_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[48]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n396), .QN(n1290) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_47_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[47]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .Q(n397), .QN(n1289) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_46_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[46]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .Q(n398), .QN(n1288) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_45_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[45]), .SI(1'b0), .E(n1010), .SE(1'b0), 
        .CK(clk), .Q(n399), .QN(n1287) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_44_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[44]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n400), .QN(n1286) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_43_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[43]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .Q(n401), .QN(n1285) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_42_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[42]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n402), .QN(n1284) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_41_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[41]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n403), .QN(n1283) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_40_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[40]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .Q(n404), .QN(n1282) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_39_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[39]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .Q(n411), .QN(n1281) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_38_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[38]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .Q(n412), .QN(n1280) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_37_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[37]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n413), .QN(n1279) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_36_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[36]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .Q(n405), .QN(n1278) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_35_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[35]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .Q(n414), .QN(n1277) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_34_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[34]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n415), .QN(n1276) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_33_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[33]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n416), .QN(n1275) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_32_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[32]), .SI(1'b0), .E(n1005), .SE(1'b0), 
        .CK(clk), .Q(n417), .QN(n1274) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_31_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[31]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .Q(n418), .QN(n1273) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_30_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[30]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n419), .QN(n1272) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_29_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[29]), .SI(1'b0), .E(n1020), .SE(1'b0), 
        .CK(clk), .Q(n420), .QN(n1271) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_28_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[28]), .SI(1'b0), .E(n1015), .SE(1'b0), 
        .CK(clk), .Q(n421), .QN(n1270) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_27_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[27]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .Q(n422), .QN(n1269) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_26_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[26]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .Q(n423), .QN(n1268) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_25_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[25]), .SI(1'b0), .E(n1014), .SE(1'b0), 
        .CK(clk), .Q(n424), .QN(n1267) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_24_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[24]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .Q(n425), .QN(n1266) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_23_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[23]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .Q(n426), .QN(n1265) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_22_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[22]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .Q(n427), .QN(n1264) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_21_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[21]), .SI(1'b0), .E(n1013), .SE(1'b0), 
        .CK(clk), .Q(n428), .QN(n1263) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_20_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[20]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .Q(n339), .QN(n1262) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_19_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[19]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .Q(n340), .QN(n1261) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_18_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[18]), .SI(1'b0), .E(n1017), .SE(1'b0), 
        .CK(clk), .Q(n429), .QN(n1260) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_17_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[17]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .Q(n430), .QN(n1259) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_16_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[16]), .SI(1'b0), .E(n1006), .SE(1'b0), 
        .CK(clk), .Q(n406), .QN(n1258) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_15_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[15]), .SI(1'b0), .E(n1011), .SE(1'b0), 
        .CK(clk), .Q(n407), .QN(n1257) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_14_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[14]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n408), .QN(n1256) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_13_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[13]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .Q(n431), .QN(n1255) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_12_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[12]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .Q(n432), .QN(n1254) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_11_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[11]), .SI(1'b0), .E(n1008), .SE(1'b0), 
        .CK(clk), .Q(n433), .QN(n1253) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_10_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[10]), .SI(1'b0), .E(n1012), .SE(1'b0), 
        .CK(clk), .Q(n434), .QN(n1252) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_9_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[9]), .SI(1'b0), .E(n1023), .SE(1'b0), 
        .CK(clk), .Q(n409), .QN(n1251) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_8_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[8]), .SI(1'b0), .E(n1026), .SE(1'b0), 
        .CK(clk), .Q(n410), .QN(n1250) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_7_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[7]), .SI(1'b0), .E(n1025), .SE(1'b0), 
        .CK(clk), .QN(n1249) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_6_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[6]), .SI(1'b0), .E(n1027), .SE(1'b0), 
        .CK(clk), .QN(n1248) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_5_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[5]), .SI(1'b0), .E(n1021), .SE(1'b0), 
        .CK(clk), .QN(n1247) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_4_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[4]), .SI(1'b0), .E(n1024), .SE(1'b0), 
        .CK(clk), .QN(n1246) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_3_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[3]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1245) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_2_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[2]), .SI(1'b0), .E(n1016), .SE(1'b0), 
        .CK(clk), .QN(n1244) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_1_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[1]), .SI(1'b0), .E(n1007), .SE(1'b0), 
        .CK(clk), .QN(n1243) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_0_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[0]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .Q(n378), .QN(n1242) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_ostate_reg_64_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_istate[64]), .SI(1'b0), .E(n1004), .SE(1'b0), 
        .CK(clk), .QN(n1241) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_0_ ( .D(Inst_AEAD_bdi[0]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1240) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_1_ ( .D(Inst_AEAD_bdi[1]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1239) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_2_ ( .D(Inst_AEAD_bdi[2]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1238) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_3_ ( .D(Inst_AEAD_bdi[3]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1237) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_4_ ( .D(Inst_AEAD_bdi[4]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1236) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_5_ ( .D(Inst_AEAD_bdi[5]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1235) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_6_ ( .D(Inst_AEAD_bdi[6]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1234) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_7_ ( .D(Inst_AEAD_bdi[7]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1233) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_8_ ( .D(Inst_AEAD_bdi[8]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1232) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_9_ ( .D(Inst_AEAD_bdi[9]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1231) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_10_ ( .D(Inst_AEAD_bdi[10]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1230) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_11_ ( .D(Inst_AEAD_bdi[11]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1229) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_12_ ( .D(Inst_AEAD_bdi[12]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1228) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_13_ ( .D(Inst_AEAD_bdi[13]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1227) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_14_ ( .D(Inst_AEAD_bdi[14]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1226) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_15_ ( .D(Inst_AEAD_bdi[15]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1225) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_16_ ( .D(Inst_AEAD_bdi[16]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1224) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_17_ ( .D(Inst_AEAD_bdi[17]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1223) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_18_ ( .D(Inst_AEAD_bdi[18]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1222) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_19_ ( .D(Inst_AEAD_bdi[19]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1221) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_20_ ( .D(Inst_AEAD_bdi[20]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1220) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_21_ ( .D(Inst_AEAD_bdi[21]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1219) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_22_ ( .D(Inst_AEAD_bdi[22]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1218) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_23_ ( .D(Inst_AEAD_bdi[23]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1217) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_24_ ( .D(Inst_AEAD_bdi[24]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1216) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_25_ ( .D(Inst_AEAD_bdi[25]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1215) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_26_ ( .D(Inst_AEAD_bdi[26]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1214) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_27_ ( .D(Inst_AEAD_bdi[27]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1213) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_28_ ( .D(Inst_AEAD_bdi[28]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1212) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_29_ ( .D(Inst_AEAD_bdi[29]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1211) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_30_ ( .D(Inst_AEAD_bdi[30]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1210) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_31_ ( .D(Inst_AEAD_bdi[31]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1209) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_32_ ( .D(Inst_AEAD_bdi[32]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1208) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_33_ ( .D(Inst_AEAD_bdi[33]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1207) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_34_ ( .D(Inst_AEAD_bdi[34]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1206) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_35_ ( .D(Inst_AEAD_bdi[35]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1205) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_36_ ( .D(Inst_AEAD_bdi[36]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1204) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_37_ ( .D(Inst_AEAD_bdi[37]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1203) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_38_ ( .D(Inst_AEAD_bdi[38]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1202) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_39_ ( .D(Inst_AEAD_bdi[39]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1201) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_40_ ( .D(Inst_AEAD_bdi[40]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1200) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_41_ ( .D(Inst_AEAD_bdi[41]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1199) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_42_ ( .D(Inst_AEAD_bdi[42]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1198) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_43_ ( .D(Inst_AEAD_bdi[43]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1197) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_44_ ( .D(Inst_AEAD_bdi[44]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1196) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_45_ ( .D(Inst_AEAD_bdi[45]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1195) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_46_ ( .D(Inst_AEAD_bdi[46]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1194) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_47_ ( .D(Inst_AEAD_bdi[47]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1193) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_48_ ( .D(Inst_AEAD_bdi[48]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1192) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_49_ ( .D(Inst_AEAD_bdi[49]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1191) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_50_ ( .D(Inst_AEAD_bdi[50]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1190) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_51_ ( .D(Inst_AEAD_bdi[51]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1189) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_52_ ( .D(Inst_AEAD_bdi[52]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1188) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_53_ ( .D(Inst_AEAD_bdi[53]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1187) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_54_ ( .D(Inst_AEAD_bdi[54]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1186) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_55_ ( .D(Inst_AEAD_bdi[55]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1185) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_56_ ( .D(Inst_AEAD_bdi[56]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1184) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_57_ ( .D(Inst_AEAD_bdi[57]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1183) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_58_ ( .D(Inst_AEAD_bdi[58]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1182) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_59_ ( .D(Inst_AEAD_bdi[59]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1181) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_60_ ( .D(Inst_AEAD_bdi[60]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1180) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_61_ ( .D(Inst_AEAD_bdi[61]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1179) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_62_ ( .D(Inst_AEAD_bdi[62]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1178) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_npub_hi_reg_63_ ( .D(Inst_AEAD_bdi[63]), 
        .SI(1'b0), .E(n470), .SE(1'b0), .CK(clk), .QN(n1177) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_96_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_64_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .QN(n1176) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_97_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_65_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .QN(n1172) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_98_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_66_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .QN(n1168) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_99_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_67_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .QN(n1164) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_100_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_68_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .QN(n1160) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_101_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_69_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .QN(n1156) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_102_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_70_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .QN(n1152) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_103_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_71_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .QN(n1148) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_104_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_72_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .QN(n1144) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_105_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_73_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .QN(n1140) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_106_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_74_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .QN(n1136) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_107_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_75_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .QN(n1132) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_108_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_76_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .QN(n1128) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_109_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_77_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .QN(n1124) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_110_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_78_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .QN(n1120) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_111_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_79_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .QN(n1116) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_112_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_80_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .QN(n1112) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_113_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_81_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .QN(n1108) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_114_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_82_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .QN(n1104) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_115_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_83_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .QN(n1100) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_116_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_84_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .QN(n1096) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_117_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_85_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .QN(n1092) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_118_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_86_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .QN(n1088) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_119_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_87_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .QN(n1084) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_120_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_88_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .QN(n1080) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_121_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_89_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .QN(n1076) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_122_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_90_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .QN(n1072) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_123_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_91_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .QN(n1068) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_124_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_92_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .QN(n1064) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_125_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_93_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .QN(n1060) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_126_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_94_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .QN(n1056) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_127_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_95_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .QN(n1052) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_ctrl_is_decrypt_reg ( .D(Inst_AEAD_decrypt), 
        .SI(1'b0), .E(n5073), .SE(1'b0), .CK(clk), .Q(n442), .QN(
        Inst_AEAD_u_cc_u_cc_ctrl_n52) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_39_ ( .D(Inst_AEAD_bdi[7]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[39]), .QN(n1603) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_47_ ( .D(Inst_AEAD_bdi[15]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[47]), .QN(n1602) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_55_ ( .D(Inst_AEAD_bdi[23]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[55]), .QN(n1601) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_63_ ( .D(Inst_AEAD_bdi[31]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[63]), .QN(n1600) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_1_ ( .D(n1047), .SI(1'b0), .E(n472), 
        .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[1]) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_2_ ( .D(n1048), .SI(1'b0), .E(n472), 
        .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[2]) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_3_ ( .D(Inst_AEAD_u_input_vbytes_3_), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[3])
         );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_0_ ( .D(Inst_AEAD_u_input_n85), 
        .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_bdi_valid_bytes[0]) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_32_ ( .D(Inst_AEAD_bdi[0]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[32]), .QN(n1595) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_33_ ( .D(Inst_AEAD_bdi[1]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[33]), .QN(n1594) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_34_ ( .D(Inst_AEAD_bdi[2]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[34]), .QN(n1593) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_35_ ( .D(Inst_AEAD_bdi[3]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[35]), .QN(n1592) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_36_ ( .D(Inst_AEAD_bdi[4]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[36]), .QN(n1591) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_37_ ( .D(Inst_AEAD_bdi[5]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[37]), .QN(n1590) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_38_ ( .D(Inst_AEAD_bdi[6]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[38]), .QN(n1589) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_40_ ( .D(Inst_AEAD_bdi[8]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[40]), .QN(n1588) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_41_ ( .D(Inst_AEAD_bdi[9]), .SI(1'b0), 
        .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[41]), .QN(n1587) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_42_ ( .D(Inst_AEAD_bdi[10]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[42]), .QN(n1586) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_43_ ( .D(Inst_AEAD_bdi[11]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[43]), .QN(n1585) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_44_ ( .D(Inst_AEAD_bdi[12]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[44]), .QN(n1584) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_45_ ( .D(Inst_AEAD_bdi[13]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[45]), .QN(n1583) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_46_ ( .D(Inst_AEAD_bdi[14]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[46]), .QN(n1582) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_48_ ( .D(Inst_AEAD_bdi[16]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[48]), .QN(n1581) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_49_ ( .D(Inst_AEAD_bdi[17]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[49]), .QN(n1580) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_50_ ( .D(Inst_AEAD_bdi[18]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[50]), .QN(n1579) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_51_ ( .D(Inst_AEAD_bdi[19]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[51]), .QN(n1578) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_52_ ( .D(Inst_AEAD_bdi[20]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[52]), .QN(n1577) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_53_ ( .D(Inst_AEAD_bdi[21]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[53]), .QN(n1576) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_54_ ( .D(Inst_AEAD_bdi[22]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[54]), .QN(n1575) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_56_ ( .D(Inst_AEAD_bdi[24]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[56]), .QN(n1574) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_57_ ( .D(Inst_AEAD_bdi[25]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[57]), .QN(n1573) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_58_ ( .D(Inst_AEAD_bdi[26]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[58]), .QN(n1572) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_59_ ( .D(Inst_AEAD_bdi[27]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[59]), .QN(n1571) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_60_ ( .D(Inst_AEAD_bdi[28]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[60]), .QN(n1570) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_61_ ( .D(Inst_AEAD_bdi[29]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[61]), .QN(n1569) );
  SEDFFXL Inst_AEAD_u_input_reg_data_reg_62_ ( .D(Inst_AEAD_bdi[30]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi[62]), .QN(n1568) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_64_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_32_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_64_), .QN(n1175) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_32_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_0_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_32_), .QN(n1174) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_0_ ( .D(Inst_AEAD_key[0]), .SI(
        1'b0), .E(n997), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_0_), .QN(n1173) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_65_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_33_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_65_), .QN(n1171) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_33_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_1_), .SI(1'b0), .E(n997), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_33_), .QN(n1170) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_1_ ( .D(Inst_AEAD_key[1]), .SI(
        1'b0), .E(n997), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_1_), .QN(n1169) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_66_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_34_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_66_), .QN(n1167) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_34_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_2_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_34_), .QN(n1166) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_2_ ( .D(Inst_AEAD_key[2]), .SI(
        1'b0), .E(n996), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_2_), .QN(n1165) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_67_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_35_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_67_), .QN(n1163) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_35_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_3_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_35_), .QN(n1162) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_3_ ( .D(Inst_AEAD_key[3]), .SI(
        1'b0), .E(n996), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_3_), .QN(n1161) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_68_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_36_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_68_), .QN(n1159) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_36_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_4_), .SI(1'b0), .E(n996), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_36_), .QN(n1158) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_4_ ( .D(Inst_AEAD_key[4]), .SI(
        1'b0), .E(n996), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_4_), .QN(n1157) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_69_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_37_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_69_), .QN(n1155) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_37_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_5_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_37_), .QN(n1154) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_5_ ( .D(Inst_AEAD_key[5]), .SI(
        1'b0), .E(n995), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_5_), .QN(n1153) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_70_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_38_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_70_), .QN(n1151) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_38_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_6_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_38_), .QN(n1150) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_6_ ( .D(Inst_AEAD_key[6]), .SI(
        1'b0), .E(n995), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_6_), .QN(n1149) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_71_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_39_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_71_), .QN(n1147) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_39_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_7_), .SI(1'b0), .E(n995), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_39_), .QN(n1146) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_7_ ( .D(Inst_AEAD_key[7]), .SI(
        1'b0), .E(n995), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_7_), .QN(n1145) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_72_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_40_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_72_), .QN(n1143) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_40_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_8_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_40_), .QN(n1142) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_8_ ( .D(Inst_AEAD_key[8]), .SI(
        1'b0), .E(n994), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_8_), .QN(n1141) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_73_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_41_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_73_), .QN(n1139) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_41_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_9_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_41_), .QN(n1138) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_9_ ( .D(Inst_AEAD_key[9]), .SI(
        1'b0), .E(n994), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_9_), .QN(n1137) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_74_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_42_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_74_), .QN(n1135) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_42_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_10_), .SI(1'b0), .E(n994), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_42_), .QN(n1134) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_10_ ( .D(Inst_AEAD_key[10]), .SI(
        1'b0), .E(n994), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_10_), .QN(n1133) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_75_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_43_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_75_), .QN(n1131) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_43_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_11_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_43_), .QN(n1130) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_11_ ( .D(Inst_AEAD_key[11]), .SI(
        1'b0), .E(n993), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_11_), .QN(n1129) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_76_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_44_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_76_), .QN(n1127) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_44_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_12_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_44_), .QN(n1126) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_12_ ( .D(Inst_AEAD_key[12]), .SI(
        1'b0), .E(n993), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_12_), .QN(n1125) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_77_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_45_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_77_), .QN(n1123) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_45_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_13_), .SI(1'b0), .E(n993), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_45_), .QN(n1122) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_13_ ( .D(Inst_AEAD_key[13]), .SI(
        1'b0), .E(n993), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_13_), .QN(n1121) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_78_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_46_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_78_), .QN(n1119) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_46_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_14_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_46_), .QN(n1118) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_14_ ( .D(Inst_AEAD_key[14]), .SI(
        1'b0), .E(n992), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_14_), .QN(n1117) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_79_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_47_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_79_), .QN(n1115) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_47_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_15_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_47_), .QN(n1114) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_15_ ( .D(Inst_AEAD_key[15]), .SI(
        1'b0), .E(n992), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_15_), .QN(n1113) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_80_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_48_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_80_), .QN(n1111) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_48_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_16_), .SI(1'b0), .E(n992), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_48_), .QN(n1110) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_16_ ( .D(Inst_AEAD_key[16]), .SI(
        1'b0), .E(n992), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_16_), .QN(n1109) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_81_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_49_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_81_), .QN(n1107) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_49_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_17_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_49_), .QN(n1106) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_17_ ( .D(Inst_AEAD_key[17]), .SI(
        1'b0), .E(n991), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_17_), .QN(n1105) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_82_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_50_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_82_), .QN(n1103) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_50_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_18_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_50_), .QN(n1102) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_18_ ( .D(Inst_AEAD_key[18]), .SI(
        1'b0), .E(n991), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_18_), .QN(n1101) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_83_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_51_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_83_), .QN(n1099) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_51_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_19_), .SI(1'b0), .E(n991), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_51_), .QN(n1098) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_19_ ( .D(Inst_AEAD_key[19]), .SI(
        1'b0), .E(n991), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_19_), .QN(n1097) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_84_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_52_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_84_), .QN(n1095) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_52_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_20_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_52_), .QN(n1094) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_20_ ( .D(Inst_AEAD_key[20]), .SI(
        1'b0), .E(n990), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_20_), .QN(n1093) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_85_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_53_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_85_), .QN(n1091) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_53_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_21_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_53_), .QN(n1090) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_21_ ( .D(Inst_AEAD_key[21]), .SI(
        1'b0), .E(n990), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_21_), .QN(n1089) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_86_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_54_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_86_), .QN(n1087) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_54_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_22_), .SI(1'b0), .E(n990), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_54_), .QN(n1086) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_22_ ( .D(Inst_AEAD_key[22]), .SI(
        1'b0), .E(n990), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_22_), .QN(n1085) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_87_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_55_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_87_), .QN(n1083) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_55_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_23_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_55_), .QN(n1082) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_23_ ( .D(Inst_AEAD_key[23]), .SI(
        1'b0), .E(n989), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_23_), .QN(n1081) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_88_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_56_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_88_), .QN(n1079) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_56_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_24_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_56_), .QN(n1078) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_24_ ( .D(Inst_AEAD_key[24]), .SI(
        1'b0), .E(n989), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_24_), .QN(n1077) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_89_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_57_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_89_), .QN(n1075) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_57_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_25_), .SI(1'b0), .E(n989), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_57_), .QN(n1074) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_25_ ( .D(Inst_AEAD_key[25]), .SI(
        1'b0), .E(n989), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_25_), .QN(n1073) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_90_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_58_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_90_), .QN(n1071) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_58_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_26_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_58_), .QN(n1070) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_26_ ( .D(Inst_AEAD_key[26]), .SI(
        1'b0), .E(n988), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_26_), .QN(n1069) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_91_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_59_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_91_), .QN(n1067) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_59_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_27_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_59_), .QN(n1066) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_27_ ( .D(Inst_AEAD_key[27]), .SI(
        1'b0), .E(n988), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_27_), .QN(n1065) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_92_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_60_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_92_), .QN(n1063) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_60_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_28_), .SI(1'b0), .E(n988), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_60_), .QN(n1062) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_28_ ( .D(Inst_AEAD_key[28]), .SI(
        1'b0), .E(n988), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_28_), .QN(n1061) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_93_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_61_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_93_), .QN(n1059) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_61_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_29_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_61_), .QN(n1058) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_29_ ( .D(Inst_AEAD_key[29]), .SI(
        1'b0), .E(n987), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_29_), .QN(n1057) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_94_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_62_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_94_), .QN(n1055) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_62_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_30_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_62_), .QN(n1054) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_30_ ( .D(Inst_AEAD_key[30]), .SI(
        1'b0), .E(n987), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_30_), .QN(n1053) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_95_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_63_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_95_), .QN(n1051) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_63_ ( .D(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_31_), .SI(1'b0), .E(n987), .SE(1'b0), 
        .CK(clk), .Q(Inst_AEAD_u_cc_u_cc_dp_reg_key_63_), .QN(n1050) );
  SEDFFXL Inst_AEAD_u_cc_u_cc_dp_reg_key_reg_31_ ( .D(Inst_AEAD_key[31]), .SI(
        1'b0), .E(n987), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_cc_u_cc_dp_reg_key_31_), .QN(n1049) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__18_ ( .D(1'b0), .SI(1'b0), .E(
        n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__18_)
         );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__0_ ( .D(pdi_data[0]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__0_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__1_ ( .D(pdi_data[1]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__1_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__2_ ( .D(pdi_data[2]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__2_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__3_ ( .D(pdi_data[3]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__3_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__4_ ( .D(pdi_data[4]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__4_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__5_ ( .D(pdi_data[5]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__5_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__6_ ( .D(pdi_data[6]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__6_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__7_ ( .D(pdi_data[7]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__7_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__8_ ( .D(pdi_data[8]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__8_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__9_ ( .D(pdi_data[9]), .SI(1'b0), 
        .E(n5074), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_hdr_buffer_memory_0__9_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__10_ ( .D(pdi_data[10]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__10_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__11_ ( .D(pdi_data[11]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__11_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__12_ ( .D(pdi_data[12]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__12_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__13_ ( .D(pdi_data[13]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__13_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__14_ ( .D(pdi_data[14]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__14_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__15_ ( .D(pdi_data[15]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__15_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__16_ ( .D(pdi_data[24]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__16_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__17_ ( .D(pdi_data[25]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__17_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__19_ ( .D(pdi_data[27]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__19_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__20_ ( .D(pdi_data[28]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__20_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__21_ ( .D(pdi_data[29]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__21_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__22_ ( .D(pdi_data[30]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__22_) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_memory_reg_0__23_ ( .D(pdi_data[31]), .SI(
        1'b0), .E(n5074), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_hdr_buffer_memory_0__23_) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_5_ ( .D(
        Inst_AEAD_bdi_valid_bytes[1]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[5]) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_6_ ( .D(
        Inst_AEAD_bdi_valid_bytes[2]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[6]) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_7_ ( .D(
        Inst_AEAD_bdi_valid_bytes[3]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[7]) );
  SEDFFXL Inst_AEAD_u_input_reg_vbytes_reg_4_ ( .D(
        Inst_AEAD_bdi_valid_bytes[0]), .SI(1'b0), .E(n472), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_bdi_valid_bytes[4]) );
  SEDFFXL Inst_AEAD_u_input_sgmt_eot_reg ( .D(pdi_data[25]), .SI(1'b0), .E(
        Inst_AEAD_u_input_n554), .SE(1'b0), .CK(clk), .Q(n1565) );
  SDFFTRXL Inst_AEAD_u_hdr_buffer_rdptr_reg_1_ ( .RN(
        Inst_AEAD_u_hdr_buffer_n374), .D(n981), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .QN(n1563) );
  SDFFTRXL Inst_AEAD_u_hdr_buffer_rdptr_reg_0_ ( .RN(n5084), .D(n981), .SI(
        1'b0), .SE(1'b0), .CK(clk), .Q(n376) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__18_ ( .D(n5076), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_hdr_buffer_memory_2__18_) );
  SDFFSQXL Inst_AEAD_u_input_is_extra_reg ( .D(Inst_AEAD_u_input_n542), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_is_extra)
         );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__18_ ( .D(n5075), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_hdr_buffer_memory_1__18_) );
  SEDFFXL Inst_AEAD_u_input_reg_sel_zero_reg ( .D(n5086), .SI(1'b0), .E(
        Inst_AEAD_u_input_n421), .SE(1'b0), .CK(clk), .Q(
        Inst_AEAD_u_input_reg_sel_zero) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_ovalid_reg ( .D(Inst_AEAD_u_hdr_buffer_n435), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_cmd_rd_valid)
         );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_reg_2_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n114), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_2_) );
  SDFFSQXL Inst_AEAD_u_input_vbytes_reg_3_ ( .D(n5080), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_vbytes_3_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_reg_1_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n115), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_1_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_round_reg_2_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n120), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_round_2_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_looped_reg ( .D(Inst_AEAD_u_hdr_buffer_n431), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_hdr_buffer_looped) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_reg_3_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n113), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_3_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__0_ ( .D(
        Inst_AEAD_u_hdr_buffer_n383), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__0_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__1_ ( .D(
        Inst_AEAD_u_hdr_buffer_n384), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__1_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__2_ ( .D(
        Inst_AEAD_u_hdr_buffer_n385), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__2_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__3_ ( .D(
        Inst_AEAD_u_hdr_buffer_n386), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__3_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__4_ ( .D(
        Inst_AEAD_u_hdr_buffer_n387), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__4_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__5_ ( .D(
        Inst_AEAD_u_hdr_buffer_n388), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__5_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__6_ ( .D(
        Inst_AEAD_u_hdr_buffer_n389), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__6_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__7_ ( .D(
        Inst_AEAD_u_hdr_buffer_n390), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__7_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__8_ ( .D(
        Inst_AEAD_u_hdr_buffer_n391), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__8_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__9_ ( .D(
        Inst_AEAD_u_hdr_buffer_n392), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__9_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__10_ ( .D(
        Inst_AEAD_u_hdr_buffer_n393), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__10_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__11_ ( .D(
        Inst_AEAD_u_hdr_buffer_n394), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__11_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__12_ ( .D(
        Inst_AEAD_u_hdr_buffer_n395), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__12_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__13_ ( .D(
        Inst_AEAD_u_hdr_buffer_n396), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__13_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__14_ ( .D(
        Inst_AEAD_u_hdr_buffer_n397), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__14_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__15_ ( .D(
        Inst_AEAD_u_hdr_buffer_n398), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__15_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__16_ ( .D(
        Inst_AEAD_u_hdr_buffer_n399), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__16_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__17_ ( .D(
        Inst_AEAD_u_hdr_buffer_n400), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__17_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__19_ ( .D(
        Inst_AEAD_u_hdr_buffer_n402), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__19_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__20_ ( .D(
        Inst_AEAD_u_hdr_buffer_n403), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__20_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__21_ ( .D(
        Inst_AEAD_u_hdr_buffer_n404), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__21_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__22_ ( .D(
        Inst_AEAD_u_hdr_buffer_n405), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__22_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_1__23_ ( .D(
        Inst_AEAD_u_hdr_buffer_n406), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_1__23_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__0_ ( .D(
        Inst_AEAD_u_hdr_buffer_n407), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__0_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__1_ ( .D(
        Inst_AEAD_u_hdr_buffer_n408), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__1_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__2_ ( .D(
        Inst_AEAD_u_hdr_buffer_n409), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__2_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__3_ ( .D(
        Inst_AEAD_u_hdr_buffer_n410), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__3_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__4_ ( .D(
        Inst_AEAD_u_hdr_buffer_n411), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__4_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__5_ ( .D(
        Inst_AEAD_u_hdr_buffer_n412), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__5_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__6_ ( .D(
        Inst_AEAD_u_hdr_buffer_n413), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__6_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__7_ ( .D(
        Inst_AEAD_u_hdr_buffer_n414), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__7_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__8_ ( .D(
        Inst_AEAD_u_hdr_buffer_n415), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__8_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__9_ ( .D(
        Inst_AEAD_u_hdr_buffer_n416), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__9_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__10_ ( .D(
        Inst_AEAD_u_hdr_buffer_n417), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__10_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__11_ ( .D(
        Inst_AEAD_u_hdr_buffer_n418), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__11_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__12_ ( .D(
        Inst_AEAD_u_hdr_buffer_n419), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__12_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__13_ ( .D(
        Inst_AEAD_u_hdr_buffer_n420), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__13_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__14_ ( .D(
        Inst_AEAD_u_hdr_buffer_n421), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__14_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__15_ ( .D(
        Inst_AEAD_u_hdr_buffer_n422), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__15_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__16_ ( .D(
        Inst_AEAD_u_hdr_buffer_n423), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__16_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__17_ ( .D(
        Inst_AEAD_u_hdr_buffer_n424), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__17_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__19_ ( .D(
        Inst_AEAD_u_hdr_buffer_n426), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__19_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__20_ ( .D(
        Inst_AEAD_u_hdr_buffer_n427), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__20_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__21_ ( .D(
        Inst_AEAD_u_hdr_buffer_n428), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__21_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__22_ ( .D(
        Inst_AEAD_u_hdr_buffer_n429), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__22_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_memory_reg_2__23_ ( .D(
        Inst_AEAD_u_hdr_buffer_n430), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_memory_2__23_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_is_init_dat_reg ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n116), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_is_init_dat) );
  SDFFSQXL Inst_AEAD_u_input_bdi_eot_reg ( .D(Inst_AEAD_u_input_n477), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_eot) );
  SDFFSQXL Inst_AEAD_u_input_ploc_reg_0_ ( .D(Inst_AEAD_u_input_n491), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ploc_0_)
         );
  SDFFSQXL Inst_AEAD_u_input_ploc_reg_1_ ( .D(Inst_AEAD_u_input_n490), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ploc_1_)
         );
  SDFFSQXL Inst_AEAD_u_input_req_pad_reg ( .D(Inst_AEAD_u_input_n492), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_req_pad)
         );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_7_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2199), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_7_) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_16_ ( .D(Inst_AEAD_u_input_n506), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[16]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_17_ ( .D(Inst_AEAD_u_input_n505), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[17]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_18_ ( .D(Inst_AEAD_u_input_n504), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[18]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_19_ ( .D(Inst_AEAD_u_input_n503), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[19]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_20_ ( .D(Inst_AEAD_u_input_n502), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[20]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_21_ ( .D(Inst_AEAD_u_input_n501), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[21]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_22_ ( .D(Inst_AEAD_u_input_n500), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[22]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_24_ ( .D(Inst_AEAD_u_input_n499), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[24]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_26_ ( .D(Inst_AEAD_u_input_n497), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[26]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_27_ ( .D(Inst_AEAD_u_input_n496), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[27]) );
  SDFFSQXL Inst_AEAD_u_input_reg_key_update_reg ( .D(Inst_AEAD_u_input_n522), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_key_update) );
  SDFFRQX2 Inst_REgIDst_do_reg_0_ ( .D(n5088), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n974), .Q(IDstReg[0]) );
  SDFFRQX2 Inst_REgIDst_do_reg_1_ ( .D(n5090), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n974), .Q(IDstReg[1]) );
  SDFFRQX2 Inst_REgIDst_do_reg_2_ ( .D(n5092), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n974), .Q(IDstReg[2]) );
  SDFFRQX2 Inst_REgIDst_do_reg_3_ ( .D(n5094), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n974), .Q(IDstReg[3]) );
  SDFFRQX2 Inst_REgIDst_do_reg_4_ ( .D(n5096), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[4]) );
  SDFFRQX2 Inst_REgIDst_do_reg_5_ ( .D(n5098), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[5]) );
  SDFFRQX2 Inst_REgIDst_do_reg_6_ ( .D(n5100), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[6]) );
  SDFFRQX2 Inst_REgIDst_do_reg_7_ ( .D(n5102), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[7]) );
  SDFFRQX2 Inst_REgIDst_do_reg_8_ ( .D(n5104), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[8]) );
  SDFFRQX2 Inst_REgIDst_do_reg_9_ ( .D(n5106), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[9]) );
  SDFFRQX2 Inst_REgIDst_do_reg_10_ ( .D(n5108), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[10]) );
  SDFFRQX2 Inst_REgIDst_do_reg_11_ ( .D(n5110), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[11]) );
  SDFFRQX2 Inst_REgIDst_do_reg_12_ ( .D(n5112), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[12]) );
  SDFFRQX2 Inst_REgIDst_do_reg_13_ ( .D(n5114), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[13]) );
  SDFFRQX2 Inst_REgIDst_do_reg_14_ ( .D(n5116), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[14]) );
  SDFFRQX2 Inst_REgIDst_do_reg_15_ ( .D(n5118), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n973), .Q(IDstReg[15]) );
  SDFFRQX2 Inst_REgIDst_do_reg_16_ ( .D(n5120), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[16]) );
  SDFFRQX2 Inst_REgIDst_do_reg_17_ ( .D(n5122), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[17]) );
  SDFFRQX2 Inst_REgIDst_do_reg_18_ ( .D(n5124), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[18]) );
  SDFFRQX2 Inst_REgIDst_do_reg_19_ ( .D(n5126), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[19]) );
  SDFFRQX2 Inst_REgIDst_do_reg_20_ ( .D(n5128), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[20]) );
  SDFFRQX2 Inst_REgIDst_do_reg_21_ ( .D(n5130), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[21]) );
  SDFFRQX2 Inst_REgIDst_do_reg_22_ ( .D(n5132), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[22]) );
  SDFFRQX2 Inst_REgIDst_do_reg_23_ ( .D(n5134), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[23]) );
  SDFFRQX2 Inst_REgIDst_do_reg_24_ ( .D(n5136), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[24]) );
  SDFFRQX2 Inst_REgIDst_do_reg_25_ ( .D(n5138), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[25]) );
  SDFFRQX2 Inst_REgIDst_do_reg_26_ ( .D(n5140), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[26]) );
  SDFFRQX2 Inst_REgIDst_do_reg_27_ ( .D(n5142), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n972), .Q(IDstReg[27]) );
  SDFFRQX2 Inst_REgIDst_do_reg_28_ ( .D(n5144), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[28]) );
  SDFFRQX2 Inst_REgIDst_do_reg_29_ ( .D(n5146), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[29]) );
  SDFFRQX2 Inst_REgIDst_do_reg_30_ ( .D(n5148), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[30]) );
  SDFFRQX2 Inst_REgIDst_do_reg_31_ ( .D(n5150), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[31]) );
  SDFFRQX2 Inst_REgIDst_do_reg_32_ ( .D(n5152), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[32]) );
  SDFFRQX2 Inst_REgIDst_do_reg_33_ ( .D(n5154), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[33]) );
  SDFFRQX2 Inst_REgIDst_do_reg_34_ ( .D(n5156), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[34]) );
  SDFFRQX2 Inst_REgIDst_do_reg_35_ ( .D(n5158), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[35]) );
  SDFFRQX2 Inst_REgIDst_do_reg_36_ ( .D(n5160), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[36]) );
  SDFFRQX2 Inst_REgIDst_do_reg_37_ ( .D(n5162), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[37]) );
  SDFFRQX2 Inst_REgIDst_do_reg_38_ ( .D(n5164), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[38]) );
  SDFFRQX2 Inst_REgIDst_do_reg_39_ ( .D(n5166), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n971), .Q(IDstReg[39]) );
  SDFFRQX2 Inst_REgIDst_do_reg_40_ ( .D(n5168), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[40]) );
  SDFFRQX2 Inst_REgIDst_do_reg_41_ ( .D(n5170), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[41]) );
  SDFFRQX2 Inst_REgIDst_do_reg_42_ ( .D(n5172), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[42]) );
  SDFFRQX2 Inst_REgIDst_do_reg_43_ ( .D(n5174), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[43]) );
  SDFFRQX2 Inst_REgIDst_do_reg_44_ ( .D(n5176), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[44]) );
  SDFFRQX2 Inst_REgIDst_do_reg_45_ ( .D(n5178), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[45]) );
  SDFFRQX2 Inst_REgIDst_do_reg_46_ ( .D(n5180), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[46]) );
  SDFFRQX2 Inst_REgIDst_do_reg_47_ ( .D(n5182), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[47]) );
  SDFFRQX2 Inst_REgIDst_do_reg_48_ ( .D(n5184), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[48]) );
  SDFFRQX2 Inst_REgIDst_do_reg_49_ ( .D(n5186), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[49]) );
  SDFFRQX2 Inst_REgIDst_do_reg_50_ ( .D(n5188), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[50]) );
  SDFFRQX2 Inst_REgIDst_do_reg_51_ ( .D(n5190), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n970), .Q(IDstReg[51]) );
  SDFFRQX2 Inst_REgIDst_do_reg_52_ ( .D(n5192), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[52]) );
  SDFFRQX2 Inst_REgIDst_do_reg_53_ ( .D(n5194), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[53]) );
  SDFFRQX2 Inst_REgIDst_do_reg_54_ ( .D(n5196), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[54]) );
  SDFFRQX2 Inst_REgIDst_do_reg_55_ ( .D(n5198), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[55]) );
  SDFFRQX2 Inst_REgIDst_do_reg_56_ ( .D(n5200), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[56]) );
  SDFFRQX2 Inst_REgIDst_do_reg_57_ ( .D(n5202), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[57]) );
  SDFFRQX2 Inst_REgIDst_do_reg_58_ ( .D(n5204), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[58]) );
  SDFFRQX2 Inst_REgIDst_do_reg_59_ ( .D(n5206), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[59]) );
  SDFFRQX2 Inst_REgIDst_do_reg_60_ ( .D(n5208), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[60]) );
  SDFFRQX2 Inst_REgIDst_do_reg_61_ ( .D(n5210), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[61]) );
  SDFFRQX2 Inst_REgIDst_do_reg_62_ ( .D(n5212), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[62]) );
  SDFFRQX2 Inst_REgIDst_do_reg_63_ ( .D(n5214), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n969), .Q(IDstReg[63]) );
  SDFFSQXL Inst_AEAD_u_input_ctr_reg_0_ ( .D(Inst_AEAD_u_input_n543), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ctr_0_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_4_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2202), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_4_) );
  SDFFSQXL Inst_AEAD_u_input_size_reg_1_ ( .D(Inst_AEAD_u_input_n482), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_size_1_)
         );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_7_ ( .D(n5079), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[7]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_15_ ( .D(n5078), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[15]) );
  SDFFSQXL Inst_AEAD_u_input_reg_data_reg_23_ ( .D(Inst_AEAD_u_input_n488), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[23]) );
  SDFFSQXL Inst_AEAD_u_input_size_reg_0_ ( .D(Inst_AEAD_u_input_n483), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_size_0_)
         );
  SDFFSQXL Inst_AEAD_u_input_reg_size_reg_3_ ( .D(Inst_AEAD_u_input_n478), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_size[3])
         );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_15_ ( .D(Inst_AEAD_u_input_n540), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_15_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_iready_reg ( .D(Inst_AEAD_u_hdr_buffer_n432), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_cmd_wr_ready)
         );
  SDFFSQXL Inst_AEAD_u_input_slen_reg_6_ ( .D(Inst_AEAD_u_input_n551), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_6_)
         );
  SDFFSQXL Inst_counter_counter_up_reg_63_ ( .D(Inst_counter_n132), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[63]) );
  SDFFSQXL Inst_AEAD_u_input_reg_bdi_valid_reg ( .D(Inst_AEAD_u_input_n521), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_valid) );
  SDFFSQXL Inst_AEAD_u_input_ss_reg_1_ ( .D(Inst_AEAD_u_input_n550), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ss_1_) );
  SDFFSQXL Inst_AEAD_u_input_ps_reg_0_ ( .D(Inst_AEAD_u_input_n524), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ps_0_) );
  SDFFSQXL Inst_AEAD_u_input_ps_reg_1_ ( .D(Inst_AEAD_u_input_n523), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ps_1_) );
  SDFFRQX2 Inst_RegIDt_do_reg_0_ ( .D(Inst_RegIDt_n3), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[0]) );
  SDFFRQX2 Inst_RegIDt_do_reg_1_ ( .D(Inst_RegIDt_n5), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[1]) );
  SDFFRQX2 Inst_RegIDt_do_reg_2_ ( .D(Inst_RegIDt_n7), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[2]) );
  SDFFRQX2 Inst_RegIDt_do_reg_3_ ( .D(Inst_RegIDt_n9), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[3]) );
  SDFFRQX2 Inst_RegIDt_do_reg_4_ ( .D(Inst_RegIDt_n11), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[4]) );
  SDFFRQX2 Inst_RegIDt_do_reg_5_ ( .D(Inst_RegIDt_n13), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[5]) );
  SDFFRQX2 Inst_RegIDt_do_reg_6_ ( .D(Inst_RegIDt_n15), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[6]) );
  SDFFRQX2 Inst_RegIDt_do_reg_7_ ( .D(Inst_RegIDt_n17), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n979), .Q(IDtReg[7]) );
  SDFFRQX2 Inst_RegIDt_do_reg_8_ ( .D(Inst_RegIDt_n19), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[8]) );
  SDFFRQX2 Inst_RegIDt_do_reg_9_ ( .D(Inst_RegIDt_n21), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[9]) );
  SDFFRQX2 Inst_RegIDt_do_reg_10_ ( .D(Inst_RegIDt_n23), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[10]) );
  SDFFRQX2 Inst_RegIDt_do_reg_11_ ( .D(Inst_RegIDt_n25), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[11]) );
  SDFFRQX2 Inst_RegIDt_do_reg_12_ ( .D(Inst_RegIDt_n27), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[12]) );
  SDFFRQX2 Inst_RegIDt_do_reg_13_ ( .D(Inst_RegIDt_n29), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[13]) );
  SDFFRQX2 Inst_RegIDt_do_reg_14_ ( .D(Inst_RegIDt_n31), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[14]) );
  SDFFRQX2 Inst_RegIDt_do_reg_15_ ( .D(Inst_RegIDt_n33), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[15]) );
  SDFFRQX2 Inst_RegIDt_do_reg_16_ ( .D(Inst_RegIDt_n35), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[16]) );
  SDFFRQX2 Inst_RegIDt_do_reg_17_ ( .D(Inst_RegIDt_n37), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[17]) );
  SDFFRQX2 Inst_RegIDt_do_reg_18_ ( .D(Inst_RegIDt_n39), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[18]) );
  SDFFRQX2 Inst_RegIDt_do_reg_19_ ( .D(Inst_RegIDt_n41), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n978), .Q(IDtReg[19]) );
  SDFFRQX2 Inst_RegIDt_do_reg_20_ ( .D(Inst_RegIDt_n43), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[20]) );
  SDFFRQX2 Inst_RegIDt_do_reg_21_ ( .D(Inst_RegIDt_n45), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[21]) );
  SDFFRQX2 Inst_RegIDt_do_reg_22_ ( .D(Inst_RegIDt_n47), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[22]) );
  SDFFRQX2 Inst_RegIDt_do_reg_23_ ( .D(Inst_RegIDt_n49), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[23]) );
  SDFFRQX2 Inst_RegIDt_do_reg_24_ ( .D(Inst_RegIDt_n51), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[24]) );
  SDFFRQX2 Inst_RegIDt_do_reg_25_ ( .D(Inst_RegIDt_n53), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[25]) );
  SDFFRQX2 Inst_RegIDt_do_reg_26_ ( .D(Inst_RegIDt_n55), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[26]) );
  SDFFRQX2 Inst_RegIDt_do_reg_27_ ( .D(Inst_RegIDt_n57), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[27]) );
  SDFFRQX2 Inst_RegIDt_do_reg_28_ ( .D(Inst_RegIDt_n59), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[28]) );
  SDFFRQX2 Inst_RegIDt_do_reg_29_ ( .D(Inst_RegIDt_n61), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[29]) );
  SDFFRQX2 Inst_RegIDt_do_reg_30_ ( .D(Inst_RegIDt_n63), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[30]) );
  SDFFRQX2 Inst_RegIDt_do_reg_31_ ( .D(Inst_RegIDt_n65), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n977), .Q(IDtReg[31]) );
  SDFFRQX2 Inst_RegIDt_do_reg_32_ ( .D(Inst_RegIDt_n67), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[32]) );
  SDFFRQX2 Inst_RegIDt_do_reg_33_ ( .D(Inst_RegIDt_n69), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[33]) );
  SDFFRQX2 Inst_RegIDt_do_reg_34_ ( .D(Inst_RegIDt_n71), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[34]) );
  SDFFRQX2 Inst_RegIDt_do_reg_35_ ( .D(Inst_RegIDt_n73), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[35]) );
  SDFFRQX2 Inst_RegIDt_do_reg_36_ ( .D(Inst_RegIDt_n75), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[36]) );
  SDFFRQX2 Inst_RegIDt_do_reg_37_ ( .D(Inst_RegIDt_n77), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[37]) );
  SDFFRQX2 Inst_RegIDt_do_reg_38_ ( .D(Inst_RegIDt_n79), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[38]) );
  SDFFRQX2 Inst_RegIDt_do_reg_39_ ( .D(Inst_RegIDt_n81), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[39]) );
  SDFFRQX2 Inst_RegIDt_do_reg_40_ ( .D(Inst_RegIDt_n83), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[40]) );
  SDFFRQX2 Inst_RegIDt_do_reg_41_ ( .D(Inst_RegIDt_n85), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[41]) );
  SDFFRQX2 Inst_RegIDt_do_reg_42_ ( .D(Inst_RegIDt_n87), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[42]) );
  SDFFRQX2 Inst_RegIDt_do_reg_43_ ( .D(Inst_RegIDt_n89), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n976), .Q(IDtReg[43]) );
  SDFFRQX2 Inst_RegIDt_do_reg_44_ ( .D(Inst_RegIDt_n91), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[44]) );
  SDFFRQX2 Inst_RegIDt_do_reg_45_ ( .D(Inst_RegIDt_n93), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[45]) );
  SDFFRQX2 Inst_RegIDt_do_reg_46_ ( .D(Inst_RegIDt_n95), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[46]) );
  SDFFRQX2 Inst_RegIDt_do_reg_47_ ( .D(Inst_RegIDt_n97), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[47]) );
  SDFFRQX2 Inst_RegIDt_do_reg_48_ ( .D(Inst_RegIDt_n99), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[48]) );
  SDFFRQX2 Inst_RegIDt_do_reg_49_ ( .D(Inst_RegIDt_n101), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[49]) );
  SDFFRQX2 Inst_RegIDt_do_reg_50_ ( .D(Inst_RegIDt_n103), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[50]) );
  SDFFRQX2 Inst_RegIDt_do_reg_51_ ( .D(Inst_RegIDt_n105), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[51]) );
  SDFFRQX2 Inst_RegIDt_do_reg_52_ ( .D(Inst_RegIDt_n107), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[52]) );
  SDFFRQX2 Inst_RegIDt_do_reg_53_ ( .D(Inst_RegIDt_n109), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[53]) );
  SDFFRQX2 Inst_RegIDt_do_reg_54_ ( .D(Inst_RegIDt_n111), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[54]) );
  SDFFRQX2 Inst_RegIDt_do_reg_55_ ( .D(Inst_RegIDt_n113), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n975), .Q(IDtReg[55]) );
  SDFFRQX2 Inst_RegIDt_do_reg_56_ ( .D(Inst_RegIDt_n115), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[56]) );
  SDFFRQX2 Inst_RegIDt_do_reg_57_ ( .D(Inst_RegIDt_n117), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[57]) );
  SDFFRQX2 Inst_RegIDt_do_reg_58_ ( .D(Inst_RegIDt_n119), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[58]) );
  SDFFRQX2 Inst_RegIDt_do_reg_59_ ( .D(Inst_RegIDt_n121), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[59]) );
  SDFFRQX2 Inst_RegIDt_do_reg_60_ ( .D(Inst_RegIDt_n123), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[60]) );
  SDFFRQX2 Inst_RegIDt_do_reg_61_ ( .D(Inst_RegIDt_n125), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[61]) );
  SDFFRQX2 Inst_RegIDt_do_reg_62_ ( .D(Inst_RegIDt_n127), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[62]) );
  SDFFRQX2 Inst_RegIDt_do_reg_63_ ( .D(Inst_RegIDt_n130), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n974), .Q(IDtReg[63]) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_0_ ( .D(Inst_AEAD_u_input_n539), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_N128)
         );
  SDFFSQXL Inst_AEAD_u_input_reg_size_reg_0_ ( .D(Inst_AEAD_u_input_n481), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_size[0])
         );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_wrptr_reg_0_ ( .D(
        Inst_AEAD_u_hdr_buffer_n433), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_wrptr_0_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_2_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2204), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_2_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_0_ ( .D(n5083), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_cc_u_cc_dp_rc_0_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_5_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2201), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_5_) );
  SDFFSX2 Inst_AEAD_u_input_slen_reg_0_ ( .D(Inst_AEAD_u_input_n552), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .QN(Inst_AEAD_u_input_n362) );
  SDFFSX2 Inst_AEAD_u_cc_u_cc_ctrl_round_reg_3_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n123), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .QN(Inst_AEAD_u_cc_u_cc_ctrl_n37) );
  SDFFSQXL Inst_AEAD_u_input_reg_size_reg_1_ ( .D(Inst_AEAD_u_input_n480), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_size[1])
         );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_state_reg_0_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n118), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_state_0_) );
  SDFFSQXL Inst_AEAD_u_input_ps_reg_2_ ( .D(Inst_AEAD_u_input_n541), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ps_2_) );
  SDFFSQXL Inst_AEAD_u_hdr_buffer_wrptr_reg_1_ ( .D(
        Inst_AEAD_u_hdr_buffer_n434), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_hdr_buffer_wrptr_1_) );
  SDFFSX2 Inst_AEAD_u_input_vbytes_reg_1_ ( .D(Inst_AEAD_u_input_n485), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(n1047), .QN(
        Inst_AEAD_u_input_n287) );
  SDFFSX2 Inst_AEAD_u_input_vbytes_reg_2_ ( .D(Inst_AEAD_u_input_n484), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(n1048), .QN(
        Inst_AEAD_u_input_n286) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_1_ ( .D(Inst_AEAD_u_input_n538), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_1_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_dp_rc_reg_1_ ( .D(n5082), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_cc_u_cc_dp_rc_1_) );
  SDFFSQXL Inst_AEAD_u_input_reg_size_reg_2_ ( .D(Inst_AEAD_u_input_n479), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi_size[2])
         );
  SDFFSX2 Inst_AEAD_u_input_ploc_reg_3_ ( .D(Inst_AEAD_u_input_n487), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .QN(n467) );
  SDFFSX2 Inst_AEAD_u_input_slen_reg_1_ ( .D(Inst_AEAD_u_input_n548), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_1_), .QN(n466) );
  SDFFSX2 Inst_AEAD_u_cc_u_cc_dp_rc_reg_6_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2200), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_6_), .QN(n377) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_state_reg_1_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n117), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_state_1_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_state_reg_2_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n119), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_state_2_) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_31_ ( .D(Inst_AEAD_u_input_n486), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[31]), .QN(
        Inst_AEAD_u_input_n303) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_0_ ( .D(Inst_AEAD_u_input_n520), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[0]), .QN(
        Inst_AEAD_u_input_n321) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_1_ ( .D(Inst_AEAD_u_input_n519), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[1]), .QN(
        Inst_AEAD_u_input_n320) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_2_ ( .D(Inst_AEAD_u_input_n518), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[2]), .QN(
        Inst_AEAD_u_input_n319) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_3_ ( .D(Inst_AEAD_u_input_n517), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[3]), .QN(
        Inst_AEAD_u_input_n318) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_4_ ( .D(Inst_AEAD_u_input_n516), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[4]), .QN(
        Inst_AEAD_u_input_n317) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_5_ ( .D(Inst_AEAD_u_input_n515), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[5]), .QN(
        Inst_AEAD_u_input_n316) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_6_ ( .D(Inst_AEAD_u_input_n514), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[6]), .QN(
        Inst_AEAD_u_input_n315) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_8_ ( .D(Inst_AEAD_u_input_n513), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[8]), .QN(
        Inst_AEAD_u_input_n314) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_9_ ( .D(Inst_AEAD_u_input_n512), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[9]), .QN(
        Inst_AEAD_u_input_n313) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_10_ ( .D(Inst_AEAD_u_input_n511), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[10]), .QN(
        Inst_AEAD_u_input_n312) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_11_ ( .D(Inst_AEAD_u_input_n510), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[11]), .QN(
        Inst_AEAD_u_input_n311) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_12_ ( .D(Inst_AEAD_u_input_n509), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[12]), .QN(
        Inst_AEAD_u_input_n310) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_13_ ( .D(Inst_AEAD_u_input_n508), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[13]), .QN(
        Inst_AEAD_u_input_n309) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_14_ ( .D(Inst_AEAD_u_input_n507), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[14]), .QN(
        Inst_AEAD_u_input_n308) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_25_ ( .D(Inst_AEAD_u_input_n498), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[25]), .QN(
        Inst_AEAD_u_input_n307) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_28_ ( .D(Inst_AEAD_u_input_n495), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[28]), .QN(
        Inst_AEAD_u_input_n306) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_29_ ( .D(Inst_AEAD_u_input_n494), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[29]), .QN(
        Inst_AEAD_u_input_n305) );
  SDFFSX2 Inst_AEAD_u_input_reg_data_reg_30_ ( .D(Inst_AEAD_u_input_n493), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_bdi[30]), .QN(
        Inst_AEAD_u_input_n304) );
  SDFFSQXL Inst_counter_counter_up_reg_0_ ( .D(Inst_counter_n195), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[0]) );
  SDFFSX2 Inst_AEAD_u_input_ploc_reg_2_ ( .D(Inst_AEAD_u_input_n489), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(n1045), .QN(n469) );
  SDFFSQXL Inst_AEAD_u_input_ss_reg_0_ ( .D(Inst_AEAD_u_input_n549), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_ss_0_) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_round_reg_0_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n122), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_sel_tag[0]) );
  SDFFSQXL Inst_AEAD_u_cc_u_cc_ctrl_round_reg_1_ ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n121), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_u_cc_ctrl_round_1_) );
  SDFFSX2 Inst_AEAD_u_cc_u_cc_dp_rc_reg_3_ ( .D(Inst_AEAD_u_cc_u_cc_dp_n2203), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_cc_u_cc_dp_rc_3_) );
  SDFFSQXL Inst_counter_counter_up_reg_62_ ( .D(Inst_counter_n133), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[62]) );
  SDFFSQXL Inst_counter_counter_up_reg_61_ ( .D(Inst_counter_n134), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[61]) );
  SDFFSQXL Inst_counter_counter_up_reg_60_ ( .D(Inst_counter_n135), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[60]) );
  SDFFSQXL Inst_counter_counter_up_reg_59_ ( .D(Inst_counter_n136), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[59]) );
  SDFFSQXL Inst_counter_counter_up_reg_58_ ( .D(Inst_counter_n137), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[58]) );
  SDFFSQXL Inst_counter_counter_up_reg_57_ ( .D(Inst_counter_n138), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[57]) );
  SDFFSQXL Inst_counter_counter_up_reg_56_ ( .D(Inst_counter_n139), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[56]) );
  SDFFSQXL Inst_counter_counter_up_reg_55_ ( .D(Inst_counter_n140), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[55]) );
  SDFFSQXL Inst_counter_counter_up_reg_54_ ( .D(Inst_counter_n141), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[54]) );
  SDFFSQXL Inst_counter_counter_up_reg_53_ ( .D(Inst_counter_n142), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[53]) );
  SDFFSQXL Inst_counter_counter_up_reg_52_ ( .D(Inst_counter_n143), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[52]) );
  SDFFSQXL Inst_counter_counter_up_reg_51_ ( .D(Inst_counter_n144), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[51]) );
  SDFFSQXL Inst_counter_counter_up_reg_50_ ( .D(Inst_counter_n145), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[50]) );
  SDFFSQXL Inst_counter_counter_up_reg_49_ ( .D(Inst_counter_n146), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[49]) );
  SDFFSQXL Inst_counter_counter_up_reg_48_ ( .D(Inst_counter_n147), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[48]) );
  SDFFSQXL Inst_counter_counter_up_reg_47_ ( .D(Inst_counter_n148), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[47]) );
  SDFFSQXL Inst_counter_counter_up_reg_46_ ( .D(Inst_counter_n149), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[46]) );
  SDFFSQXL Inst_counter_counter_up_reg_45_ ( .D(Inst_counter_n150), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[45]) );
  SDFFSQXL Inst_counter_counter_up_reg_44_ ( .D(Inst_counter_n151), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[44]) );
  SDFFSQXL Inst_counter_counter_up_reg_43_ ( .D(Inst_counter_n152), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[43]) );
  SDFFSQXL Inst_counter_counter_up_reg_42_ ( .D(Inst_counter_n153), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[42]) );
  SDFFSQXL Inst_counter_counter_up_reg_41_ ( .D(Inst_counter_n154), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[41]) );
  SDFFSQXL Inst_counter_counter_up_reg_40_ ( .D(Inst_counter_n155), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[40]) );
  SDFFSQXL Inst_counter_counter_up_reg_39_ ( .D(Inst_counter_n156), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[39]) );
  SDFFSQXL Inst_counter_counter_up_reg_38_ ( .D(Inst_counter_n157), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[38]) );
  SDFFSQXL Inst_counter_counter_up_reg_37_ ( .D(Inst_counter_n158), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[37]) );
  SDFFSQXL Inst_counter_counter_up_reg_36_ ( .D(Inst_counter_n159), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[36]) );
  SDFFSQXL Inst_counter_counter_up_reg_35_ ( .D(Inst_counter_n160), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[35]) );
  SDFFSQXL Inst_counter_counter_up_reg_34_ ( .D(Inst_counter_n161), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[34]) );
  SDFFSQXL Inst_counter_counter_up_reg_33_ ( .D(Inst_counter_n162), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[33]) );
  SDFFSQXL Inst_counter_counter_up_reg_32_ ( .D(Inst_counter_n163), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[32]) );
  SDFFSQXL Inst_counter_counter_up_reg_31_ ( .D(Inst_counter_n164), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[31]) );
  SDFFSQXL Inst_counter_counter_up_reg_30_ ( .D(Inst_counter_n165), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[30]) );
  SDFFSQXL Inst_counter_counter_up_reg_29_ ( .D(Inst_counter_n166), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[29]) );
  SDFFSQXL Inst_counter_counter_up_reg_28_ ( .D(Inst_counter_n167), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[28]) );
  SDFFSQXL Inst_counter_counter_up_reg_27_ ( .D(Inst_counter_n168), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[27]) );
  SDFFSQXL Inst_counter_counter_up_reg_26_ ( .D(Inst_counter_n169), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[26]) );
  SDFFSQXL Inst_counter_counter_up_reg_25_ ( .D(Inst_counter_n170), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[25]) );
  SDFFSQXL Inst_counter_counter_up_reg_24_ ( .D(Inst_counter_n171), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[24]) );
  SDFFSQXL Inst_counter_counter_up_reg_23_ ( .D(Inst_counter_n172), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[23]) );
  SDFFSQXL Inst_counter_counter_up_reg_22_ ( .D(Inst_counter_n173), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[22]) );
  SDFFSQXL Inst_counter_counter_up_reg_21_ ( .D(Inst_counter_n174), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[21]) );
  SDFFSQXL Inst_counter_counter_up_reg_20_ ( .D(Inst_counter_n175), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[20]) );
  SDFFSQXL Inst_counter_counter_up_reg_19_ ( .D(Inst_counter_n176), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[19]) );
  SDFFSQXL Inst_counter_counter_up_reg_18_ ( .D(Inst_counter_n177), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[18]) );
  SDFFSQXL Inst_counter_counter_up_reg_17_ ( .D(Inst_counter_n178), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[17]) );
  SDFFSQXL Inst_counter_counter_up_reg_16_ ( .D(Inst_counter_n179), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[16]) );
  SDFFSQXL Inst_counter_counter_up_reg_15_ ( .D(Inst_counter_n180), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[15]) );
  SDFFSQXL Inst_counter_counter_up_reg_14_ ( .D(Inst_counter_n181), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[14]) );
  SDFFSQXL Inst_counter_counter_up_reg_13_ ( .D(Inst_counter_n182), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[13]) );
  SDFFSQXL Inst_counter_counter_up_reg_12_ ( .D(Inst_counter_n183), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[12]) );
  SDFFSQXL Inst_counter_counter_up_reg_11_ ( .D(Inst_counter_n184), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[11]) );
  SDFFSQXL Inst_counter_counter_up_reg_10_ ( .D(Inst_counter_n185), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[10]) );
  SDFFSQXL Inst_counter_counter_up_reg_9_ ( .D(Inst_counter_n186), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[9]) );
  SDFFSQXL Inst_counter_counter_up_reg_8_ ( .D(Inst_counter_n187), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[8]) );
  SDFFSQXL Inst_counter_counter_up_reg_7_ ( .D(Inst_counter_n188), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[7]) );
  SDFFSQXL Inst_counter_counter_up_reg_6_ ( .D(Inst_counter_n189), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[6]) );
  SDFFSQXL Inst_counter_counter_up_reg_5_ ( .D(Inst_counter_n190), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[5]) );
  SDFFSQXL Inst_counter_counter_up_reg_4_ ( .D(Inst_counter_n191), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[4]) );
  SDFFSQXL Inst_counter_counter_up_reg_3_ ( .D(Inst_counter_n192), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[3]) );
  SDFFSQXL Inst_counter_counter_up_reg_2_ ( .D(Inst_counter_n193), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[2]) );
  SDFFSQXL Inst_counter_counter_up_reg_1_ ( .D(Inst_counter_n194), .SI(1'b0), 
        .SE(1'b0), .CK(clk), .SN(1'b1), .Q(randd[1]) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_13_ ( .D(Inst_AEAD_u_input_n526), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_13_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_14_ ( .D(Inst_AEAD_u_input_n525), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_14_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_11_ ( .D(Inst_AEAD_u_input_n528), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_11_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_6_ ( .D(Inst_AEAD_u_input_n533), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_6_) );
  SDFFSQXL Inst_AEAD_u_input_slen_reg_3_ ( .D(Inst_AEAD_u_input_n546), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_3_)
         );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_4_ ( .D(Inst_AEAD_u_input_n535), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_4_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_10_ ( .D(Inst_AEAD_u_input_n529), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_10_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_8_ ( .D(Inst_AEAD_u_input_n531), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_8_) );
  SDFFSQXL Inst_AEAD_u_input_slen_reg_5_ ( .D(Inst_AEAD_u_input_n544), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_5_)
         );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_12_ ( .D(Inst_AEAD_u_input_n527), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_12_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_7_ ( .D(Inst_AEAD_u_input_n532), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_7_) );
  SDFFSQXL Inst_AEAD_u_input_slen_reg_4_ ( .D(Inst_AEAD_u_input_n545), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_4_)
         );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_5_ ( .D(Inst_AEAD_u_input_n534), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_5_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_3_ ( .D(Inst_AEAD_u_input_n536), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_3_) );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_9_ ( .D(Inst_AEAD_u_input_n530), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_9_) );
  SDFFSQXL Inst_AEAD_u_input_slen_reg_2_ ( .D(Inst_AEAD_u_input_n547), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_input_slen_2_)
         );
  SDFFSQXL Inst_AEAD_u_input_sgmt_len_reg_2_ ( .D(Inst_AEAD_u_input_n537), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_AEAD_u_input_sgmt_len_2_) );
  SDFFSQX4 Inst_AEAD_u_cc_u_cc_ctrl_is_tag_reg ( .D(n5072), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(Inst_AEAD_u_cc_sel_tag[1]) );
  SDFFSQX4 Inst_AEAD_u_cc_u_cc_ctrl_sel_key_lo_reg ( .D(
        Inst_AEAD_u_cc_u_cc_ctrl_n112), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_AEAD_u_cc_sel_key_lo) );
  ADDHX1 Inst_counter_add_3021_U1_1_62 ( .A(randd[62]), .B(
        Inst_counter_add_3021_carry[62]), .CO(Inst_counter_add_3021_carry[63]), 
        .S(Inst_counter_N66) );
  ADDHX1 Inst_counter_add_3021_U1_1_61 ( .A(randd[61]), .B(
        Inst_counter_add_3021_carry[61]), .CO(Inst_counter_add_3021_carry[62]), 
        .S(Inst_counter_N65) );
  ADDHX1 Inst_counter_add_3021_U1_1_60 ( .A(randd[60]), .B(
        Inst_counter_add_3021_carry[60]), .CO(Inst_counter_add_3021_carry[61]), 
        .S(Inst_counter_N64) );
  ADDHX1 Inst_counter_add_3021_U1_1_59 ( .A(randd[59]), .B(
        Inst_counter_add_3021_carry[59]), .CO(Inst_counter_add_3021_carry[60]), 
        .S(Inst_counter_N63) );
  ADDHX1 Inst_counter_add_3021_U1_1_58 ( .A(randd[58]), .B(
        Inst_counter_add_3021_carry[58]), .CO(Inst_counter_add_3021_carry[59]), 
        .S(Inst_counter_N62) );
  ADDHX1 Inst_counter_add_3021_U1_1_57 ( .A(randd[57]), .B(
        Inst_counter_add_3021_carry[57]), .CO(Inst_counter_add_3021_carry[58]), 
        .S(Inst_counter_N61) );
  ADDHX1 Inst_counter_add_3021_U1_1_56 ( .A(randd[56]), .B(
        Inst_counter_add_3021_carry[56]), .CO(Inst_counter_add_3021_carry[57]), 
        .S(Inst_counter_N60) );
  ADDHX1 Inst_counter_add_3021_U1_1_55 ( .A(randd[55]), .B(
        Inst_counter_add_3021_carry[55]), .CO(Inst_counter_add_3021_carry[56]), 
        .S(Inst_counter_N59) );
  ADDHX1 Inst_counter_add_3021_U1_1_54 ( .A(randd[54]), .B(
        Inst_counter_add_3021_carry[54]), .CO(Inst_counter_add_3021_carry[55]), 
        .S(Inst_counter_N58) );
  ADDHX1 Inst_counter_add_3021_U1_1_53 ( .A(randd[53]), .B(
        Inst_counter_add_3021_carry[53]), .CO(Inst_counter_add_3021_carry[54]), 
        .S(Inst_counter_N57) );
  ADDHX1 Inst_counter_add_3021_U1_1_52 ( .A(randd[52]), .B(
        Inst_counter_add_3021_carry[52]), .CO(Inst_counter_add_3021_carry[53]), 
        .S(Inst_counter_N56) );
  ADDHX1 Inst_counter_add_3021_U1_1_51 ( .A(randd[51]), .B(
        Inst_counter_add_3021_carry[51]), .CO(Inst_counter_add_3021_carry[52]), 
        .S(Inst_counter_N55) );
  ADDHX1 Inst_counter_add_3021_U1_1_50 ( .A(randd[50]), .B(
        Inst_counter_add_3021_carry[50]), .CO(Inst_counter_add_3021_carry[51]), 
        .S(Inst_counter_N54) );
  ADDHX1 Inst_counter_add_3021_U1_1_49 ( .A(randd[49]), .B(
        Inst_counter_add_3021_carry[49]), .CO(Inst_counter_add_3021_carry[50]), 
        .S(Inst_counter_N53) );
  ADDHX1 Inst_counter_add_3021_U1_1_48 ( .A(randd[48]), .B(
        Inst_counter_add_3021_carry[48]), .CO(Inst_counter_add_3021_carry[49]), 
        .S(Inst_counter_N52) );
  ADDHX1 Inst_counter_add_3021_U1_1_47 ( .A(randd[47]), .B(
        Inst_counter_add_3021_carry[47]), .CO(Inst_counter_add_3021_carry[48]), 
        .S(Inst_counter_N51) );
  ADDHX1 Inst_counter_add_3021_U1_1_46 ( .A(randd[46]), .B(
        Inst_counter_add_3021_carry[46]), .CO(Inst_counter_add_3021_carry[47]), 
        .S(Inst_counter_N50) );
  ADDHX1 Inst_counter_add_3021_U1_1_45 ( .A(randd[45]), .B(
        Inst_counter_add_3021_carry[45]), .CO(Inst_counter_add_3021_carry[46]), 
        .S(Inst_counter_N49) );
  ADDHX1 Inst_counter_add_3021_U1_1_44 ( .A(randd[44]), .B(
        Inst_counter_add_3021_carry[44]), .CO(Inst_counter_add_3021_carry[45]), 
        .S(Inst_counter_N48) );
  ADDHX1 Inst_counter_add_3021_U1_1_43 ( .A(randd[43]), .B(
        Inst_counter_add_3021_carry[43]), .CO(Inst_counter_add_3021_carry[44]), 
        .S(Inst_counter_N47) );
  ADDHX1 Inst_counter_add_3021_U1_1_42 ( .A(randd[42]), .B(
        Inst_counter_add_3021_carry[42]), .CO(Inst_counter_add_3021_carry[43]), 
        .S(Inst_counter_N46) );
  ADDHX1 Inst_counter_add_3021_U1_1_41 ( .A(randd[41]), .B(
        Inst_counter_add_3021_carry[41]), .CO(Inst_counter_add_3021_carry[42]), 
        .S(Inst_counter_N45) );
  ADDHX1 Inst_counter_add_3021_U1_1_40 ( .A(randd[40]), .B(
        Inst_counter_add_3021_carry[40]), .CO(Inst_counter_add_3021_carry[41]), 
        .S(Inst_counter_N44) );
  ADDHX1 Inst_counter_add_3021_U1_1_39 ( .A(randd[39]), .B(
        Inst_counter_add_3021_carry[39]), .CO(Inst_counter_add_3021_carry[40]), 
        .S(Inst_counter_N43) );
  ADDHX1 Inst_counter_add_3021_U1_1_38 ( .A(randd[38]), .B(
        Inst_counter_add_3021_carry[38]), .CO(Inst_counter_add_3021_carry[39]), 
        .S(Inst_counter_N42) );
  ADDHX1 Inst_counter_add_3021_U1_1_37 ( .A(randd[37]), .B(
        Inst_counter_add_3021_carry[37]), .CO(Inst_counter_add_3021_carry[38]), 
        .S(Inst_counter_N41) );
  ADDHX1 Inst_counter_add_3021_U1_1_36 ( .A(randd[36]), .B(
        Inst_counter_add_3021_carry[36]), .CO(Inst_counter_add_3021_carry[37]), 
        .S(Inst_counter_N40) );
  ADDHX1 Inst_counter_add_3021_U1_1_35 ( .A(randd[35]), .B(
        Inst_counter_add_3021_carry[35]), .CO(Inst_counter_add_3021_carry[36]), 
        .S(Inst_counter_N39) );
  ADDHX1 Inst_counter_add_3021_U1_1_34 ( .A(randd[34]), .B(
        Inst_counter_add_3021_carry[34]), .CO(Inst_counter_add_3021_carry[35]), 
        .S(Inst_counter_N38) );
  ADDHX1 Inst_counter_add_3021_U1_1_33 ( .A(randd[33]), .B(
        Inst_counter_add_3021_carry[33]), .CO(Inst_counter_add_3021_carry[34]), 
        .S(Inst_counter_N37) );
  ADDHX1 Inst_counter_add_3021_U1_1_32 ( .A(randd[32]), .B(
        Inst_counter_add_3021_carry[32]), .CO(Inst_counter_add_3021_carry[33]), 
        .S(Inst_counter_N36) );
  ADDHX1 Inst_counter_add_3021_U1_1_31 ( .A(randd[31]), .B(
        Inst_counter_add_3021_carry[31]), .CO(Inst_counter_add_3021_carry[32]), 
        .S(Inst_counter_N35) );
  ADDHX1 Inst_counter_add_3021_U1_1_30 ( .A(randd[30]), .B(
        Inst_counter_add_3021_carry[30]), .CO(Inst_counter_add_3021_carry[31]), 
        .S(Inst_counter_N34) );
  ADDHX1 Inst_counter_add_3021_U1_1_29 ( .A(randd[29]), .B(
        Inst_counter_add_3021_carry[29]), .CO(Inst_counter_add_3021_carry[30]), 
        .S(Inst_counter_N33) );
  ADDHX1 Inst_counter_add_3021_U1_1_28 ( .A(randd[28]), .B(
        Inst_counter_add_3021_carry[28]), .CO(Inst_counter_add_3021_carry[29]), 
        .S(Inst_counter_N32) );
  ADDHX1 Inst_counter_add_3021_U1_1_27 ( .A(randd[27]), .B(
        Inst_counter_add_3021_carry[27]), .CO(Inst_counter_add_3021_carry[28]), 
        .S(Inst_counter_N31) );
  ADDHX1 Inst_counter_add_3021_U1_1_26 ( .A(randd[26]), .B(
        Inst_counter_add_3021_carry[26]), .CO(Inst_counter_add_3021_carry[27]), 
        .S(Inst_counter_N30) );
  ADDHX1 Inst_counter_add_3021_U1_1_25 ( .A(randd[25]), .B(
        Inst_counter_add_3021_carry[25]), .CO(Inst_counter_add_3021_carry[26]), 
        .S(Inst_counter_N29) );
  ADDHX1 Inst_counter_add_3021_U1_1_24 ( .A(randd[24]), .B(
        Inst_counter_add_3021_carry[24]), .CO(Inst_counter_add_3021_carry[25]), 
        .S(Inst_counter_N28) );
  ADDHX1 Inst_counter_add_3021_U1_1_23 ( .A(randd[23]), .B(
        Inst_counter_add_3021_carry[23]), .CO(Inst_counter_add_3021_carry[24]), 
        .S(Inst_counter_N27) );
  ADDHX1 Inst_counter_add_3021_U1_1_22 ( .A(randd[22]), .B(
        Inst_counter_add_3021_carry[22]), .CO(Inst_counter_add_3021_carry[23]), 
        .S(Inst_counter_N26) );
  ADDHX1 Inst_counter_add_3021_U1_1_21 ( .A(randd[21]), .B(
        Inst_counter_add_3021_carry[21]), .CO(Inst_counter_add_3021_carry[22]), 
        .S(Inst_counter_N25) );
  ADDHX1 Inst_counter_add_3021_U1_1_20 ( .A(randd[20]), .B(
        Inst_counter_add_3021_carry[20]), .CO(Inst_counter_add_3021_carry[21]), 
        .S(Inst_counter_N24) );
  ADDHX1 Inst_counter_add_3021_U1_1_19 ( .A(randd[19]), .B(
        Inst_counter_add_3021_carry[19]), .CO(Inst_counter_add_3021_carry[20]), 
        .S(Inst_counter_N23) );
  ADDHX1 Inst_counter_add_3021_U1_1_18 ( .A(randd[18]), .B(
        Inst_counter_add_3021_carry[18]), .CO(Inst_counter_add_3021_carry[19]), 
        .S(Inst_counter_N22) );
  ADDHX1 Inst_counter_add_3021_U1_1_17 ( .A(randd[17]), .B(
        Inst_counter_add_3021_carry[17]), .CO(Inst_counter_add_3021_carry[18]), 
        .S(Inst_counter_N21) );
  ADDHX1 Inst_counter_add_3021_U1_1_16 ( .A(randd[16]), .B(
        Inst_counter_add_3021_carry[16]), .CO(Inst_counter_add_3021_carry[17]), 
        .S(Inst_counter_N20) );
  ADDHX1 Inst_counter_add_3021_U1_1_15 ( .A(randd[15]), .B(
        Inst_counter_add_3021_carry[15]), .CO(Inst_counter_add_3021_carry[16]), 
        .S(Inst_counter_N19) );
  ADDHX1 Inst_counter_add_3021_U1_1_14 ( .A(randd[14]), .B(
        Inst_counter_add_3021_carry[14]), .CO(Inst_counter_add_3021_carry[15]), 
        .S(Inst_counter_N18) );
  ADDHX1 Inst_counter_add_3021_U1_1_13 ( .A(randd[13]), .B(
        Inst_counter_add_3021_carry[13]), .CO(Inst_counter_add_3021_carry[14]), 
        .S(Inst_counter_N17) );
  ADDHX1 Inst_counter_add_3021_U1_1_12 ( .A(randd[12]), .B(
        Inst_counter_add_3021_carry[12]), .CO(Inst_counter_add_3021_carry[13]), 
        .S(Inst_counter_N16) );
  ADDHX1 Inst_counter_add_3021_U1_1_11 ( .A(randd[11]), .B(
        Inst_counter_add_3021_carry[11]), .CO(Inst_counter_add_3021_carry[12]), 
        .S(Inst_counter_N15) );
  ADDHX1 Inst_counter_add_3021_U1_1_10 ( .A(randd[10]), .B(
        Inst_counter_add_3021_carry[10]), .CO(Inst_counter_add_3021_carry[11]), 
        .S(Inst_counter_N14) );
  ADDHX1 Inst_counter_add_3021_U1_1_9 ( .A(randd[9]), .B(
        Inst_counter_add_3021_carry[9]), .CO(Inst_counter_add_3021_carry[10]), 
        .S(Inst_counter_N13) );
  ADDHX1 Inst_counter_add_3021_U1_1_8 ( .A(randd[8]), .B(
        Inst_counter_add_3021_carry[8]), .CO(Inst_counter_add_3021_carry[9]), 
        .S(Inst_counter_N12) );
  ADDHX1 Inst_counter_add_3021_U1_1_7 ( .A(randd[7]), .B(
        Inst_counter_add_3021_carry[7]), .CO(Inst_counter_add_3021_carry[8]), 
        .S(Inst_counter_N11) );
  ADDHX1 Inst_counter_add_3021_U1_1_6 ( .A(randd[6]), .B(
        Inst_counter_add_3021_carry[6]), .CO(Inst_counter_add_3021_carry[7]), 
        .S(Inst_counter_N10) );
  ADDHX1 Inst_counter_add_3021_U1_1_5 ( .A(randd[5]), .B(
        Inst_counter_add_3021_carry[5]), .CO(Inst_counter_add_3021_carry[6]), 
        .S(Inst_counter_N9) );
  ADDHX1 Inst_counter_add_3021_U1_1_4 ( .A(randd[4]), .B(
        Inst_counter_add_3021_carry[4]), .CO(Inst_counter_add_3021_carry[5]), 
        .S(Inst_counter_N8) );
  ADDHX1 Inst_counter_add_3021_U1_1_3 ( .A(randd[3]), .B(
        Inst_counter_add_3021_carry[3]), .CO(Inst_counter_add_3021_carry[4]), 
        .S(Inst_counter_N7) );
  ADDHX1 Inst_counter_add_3021_U1_1_2 ( .A(randd[2]), .B(
        Inst_counter_add_3021_carry[2]), .CO(Inst_counter_add_3021_carry[3]), 
        .S(Inst_counter_N6) );
  ADDHX1 Inst_counter_add_3021_U1_1_1 ( .A(randd[1]), .B(randd[0]), .CO(
        Inst_counter_add_3021_carry[2]), .S(Inst_counter_N5) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_0_ ( .D(Inst_AEAD_u_hdr_buffer_N366), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[0]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_1_ ( .D(Inst_AEAD_u_hdr_buffer_N365), 
        .SI(1'b0), .E(n981), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[1]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_2_ ( .D(Inst_AEAD_u_hdr_buffer_N364), 
        .SI(1'b0), .E(n981), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[2]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_3_ ( .D(Inst_AEAD_u_hdr_buffer_N363), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[3]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_4_ ( .D(Inst_AEAD_u_hdr_buffer_N362), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[4]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_5_ ( .D(Inst_AEAD_u_hdr_buffer_N361), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[5]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_6_ ( .D(Inst_AEAD_u_hdr_buffer_N360), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[6]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_7_ ( .D(Inst_AEAD_u_hdr_buffer_N359), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[7]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_8_ ( .D(Inst_AEAD_u_hdr_buffer_N358), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[8]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_9_ ( .D(Inst_AEAD_u_hdr_buffer_N357), 
        .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[9]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_10_ ( .D(Inst_AEAD_u_hdr_buffer_N356), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[10]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_11_ ( .D(Inst_AEAD_u_hdr_buffer_N355), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[11]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_12_ ( .D(Inst_AEAD_u_hdr_buffer_N354), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[12]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_13_ ( .D(Inst_AEAD_u_hdr_buffer_N353), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[13]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_14_ ( .D(Inst_AEAD_u_hdr_buffer_N352), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[14]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_15_ ( .D(Inst_AEAD_u_hdr_buffer_N351), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[15]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_16_ ( .D(Inst_AEAD_u_hdr_buffer_N350), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[16]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_17_ ( .D(Inst_AEAD_u_hdr_buffer_N349), .SI(1'b0), .E(n980), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[17]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_18_ ( .D(Inst_AEAD_u_hdr_buffer_N348), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[18]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_19_ ( .D(Inst_AEAD_u_hdr_buffer_N347), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[19]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_20_ ( .D(Inst_AEAD_u_hdr_buffer_N346), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[20]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_21_ ( .D(Inst_AEAD_u_hdr_buffer_N345), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[21]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_22_ ( .D(Inst_AEAD_u_hdr_buffer_N344), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[22]) );
  SEDFFXL Inst_AEAD_u_hdr_buffer_dout_reg_23_ ( .D(Inst_AEAD_u_hdr_buffer_N343), .SI(1'b0), .E(n979), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_cmd_dout[23]) );
  SEDFFXL Inst_AEAD_u_input_is_decrypt_reg ( .D(pdi_data[28]), .SI(1'b0), .E(
        Inst_AEAD_u_input_n553), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_decrypt) );
  SEDFFXL Inst_AEAD_u_input_vbytes_reg_0_ ( .D(n5085), .SI(1'b0), .E(
        Inst_AEAD_u_input_n392), .SE(1'b0), .CK(clk), .Q(Inst_AEAD_u_input_n85) );
  OR2X2 U368 ( .A(n1763), .B(n2900), .Y(n337) );
  OR3X2 U369 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_0_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .C(n4367), .Y(n338) );
  NOR2X2 U370 ( .A(n1629), .B(rst), .Y(n1628) );
  NOR2X4 U371 ( .A(rst), .B(en_c), .Y(n1629) );
  NAND2BX2 U372 ( .AN(Inst_AEAD_u_cc_sel_tag[0]), .B(Inst_AEAD_u_cc_sel_tag[1]), .Y(n4931) );
  NAND3X4 U373 ( .A(n4915), .B(n4917), .C(MuxSel1[0]), .Y(n4473) );
  NAND3X4 U374 ( .A(n4915), .B(n4917), .C(n4920), .Y(n4478) );
  INVX4 U375 ( .A(n338), .Y(n470) );
  INVXL U376 ( .A(Inst_AEAD_u_input_n391), .Y(n471) );
  INVX4 U377 ( .A(n471), .Y(n472) );
  NOR3X2 U378 ( .A(Inst_AEAD_u_hdr_buffer_n374), .B(n1822), .C(n1785), .Y(
        n1796) );
  NAND3X2 U379 ( .A(MuxSel1[0]), .B(n4915), .C(MuxSel2), .Y(n4474) );
  NAND3X2 U380 ( .A(n5084), .B(n1788), .C(Inst_AEAD_u_hdr_buffer_n374), .Y(
        n1793) );
  NOR2X2 U381 ( .A(rst), .B(n1610), .Y(n5074) );
  NOR2X2 U382 ( .A(n1788), .B(rst), .Y(Inst_AEAD_u_hdr_buffer_n326) );
  NAND2X2 U383 ( .A(n1787), .B(Inst_AEAD_u_hdr_buffer_wrptr_1_), .Y(n1788) );
  NOR2X4 U384 ( .A(n1791), .B(rst), .Y(n1611) );
  NAND2XL U385 ( .A(n1787), .B(n1827), .Y(n1791) );
  NOR2X4 U386 ( .A(n1790), .B(rst), .Y(n1612) );
  NAND3X2 U387 ( .A(n4920), .B(n4915), .C(MuxSel2), .Y(n4479) );
  BUFX2 U388 ( .A(n964), .Y(n953) );
  BUFX2 U389 ( .A(n964), .Y(n954) );
  BUFX2 U390 ( .A(n964), .Y(n955) );
  BUFX2 U391 ( .A(n963), .Y(n956) );
  BUFX2 U392 ( .A(n963), .Y(n957) );
  BUFX2 U393 ( .A(n963), .Y(n958) );
  BUFX2 U394 ( .A(n966), .Y(n964) );
  BUFX2 U395 ( .A(n966), .Y(n963) );
  BUFX2 U396 ( .A(n965), .Y(n952) );
  BUFX2 U397 ( .A(n966), .Y(n965) );
  BUFX2 U398 ( .A(n962), .Y(n959) );
  BUFX2 U399 ( .A(n962), .Y(n960) );
  BUFX2 U400 ( .A(n962), .Y(n961) );
  BUFX2 U401 ( .A(n967), .Y(n962) );
  BUFX2 U402 ( .A(n968), .Y(n967) );
  BUFX2 U403 ( .A(n968), .Y(n966) );
  BUFX2 U404 ( .A(n914), .Y(n887) );
  BUFX2 U405 ( .A(n908), .Y(n906) );
  BUFX2 U406 ( .A(n913), .Y(n891) );
  BUFX2 U407 ( .A(n913), .Y(n890) );
  BUFX2 U408 ( .A(n914), .Y(n889) );
  BUFX2 U409 ( .A(n914), .Y(n888) );
  BUFX2 U410 ( .A(n913), .Y(n892) );
  BUFX2 U411 ( .A(n908), .Y(n905) );
  BUFX2 U412 ( .A(n911), .Y(n896) );
  BUFX2 U413 ( .A(n912), .Y(n895) );
  BUFX2 U414 ( .A(n912), .Y(n894) );
  BUFX2 U415 ( .A(n912), .Y(n893) );
  BUFX2 U416 ( .A(n911), .Y(n897) );
  BUFX2 U417 ( .A(n911), .Y(n898) );
  BUFX2 U418 ( .A(n910), .Y(n899) );
  BUFX2 U419 ( .A(n910), .Y(n900) );
  BUFX2 U420 ( .A(n910), .Y(n901) );
  BUFX2 U421 ( .A(n909), .Y(n902) );
  BUFX2 U422 ( .A(n909), .Y(n904) );
  BUFX2 U423 ( .A(n909), .Y(n903) );
  BUFX2 U424 ( .A(n915), .Y(n886) );
  BUFX2 U425 ( .A(n915), .Y(n885) );
  BUFX2 U426 ( .A(n915), .Y(n884) );
  INVX2 U427 ( .A(n937), .Y(n917) );
  INVX2 U428 ( .A(n942), .Y(n927) );
  INVX2 U429 ( .A(n944), .Y(n931) );
  INVX2 U430 ( .A(n944), .Y(n930) );
  INVX2 U431 ( .A(n943), .Y(n929) );
  INVX2 U432 ( .A(n943), .Y(n928) );
  INVX2 U433 ( .A(n941), .Y(n926) );
  INVX2 U434 ( .A(n941), .Y(n925) );
  INVX2 U435 ( .A(n940), .Y(n923) );
  INVX2 U436 ( .A(n939), .Y(n922) );
  INVX2 U437 ( .A(n939), .Y(n921) );
  INVX2 U438 ( .A(n942), .Y(n920) );
  INVX2 U439 ( .A(n940), .Y(n924) );
  INVX2 U440 ( .A(n938), .Y(n919) );
  INVX2 U441 ( .A(n938), .Y(n918) );
  BUFX2 U442 ( .A(n908), .Y(n907) );
  BUFX2 U443 ( .A(n1857), .Y(n910) );
  BUFX2 U444 ( .A(n1857), .Y(n908) );
  BUFX2 U445 ( .A(n1857), .Y(n909) );
  BUFX2 U446 ( .A(n1857), .Y(n911) );
  BUFX2 U447 ( .A(n1857), .Y(n912) );
  BUFX2 U448 ( .A(n1857), .Y(n913) );
  BUFX2 U449 ( .A(n1857), .Y(n914) );
  BUFX2 U450 ( .A(n1857), .Y(n915) );
  BUFX2 U451 ( .A(n951), .Y(n937) );
  BUFX2 U452 ( .A(n950), .Y(n941) );
  BUFX2 U453 ( .A(n950), .Y(n939) );
  BUFX2 U454 ( .A(n949), .Y(n944) );
  BUFX2 U455 ( .A(n949), .Y(n943) );
  BUFX2 U456 ( .A(n949), .Y(n942) );
  BUFX2 U457 ( .A(n950), .Y(n940) );
  BUFX2 U458 ( .A(n951), .Y(n938) );
  BUFX2 U459 ( .A(n2923), .Y(n968) );
  BUFX2 U460 ( .A(n1036), .Y(n1007) );
  BUFX2 U461 ( .A(n1037), .Y(n1002) );
  BUFX2 U462 ( .A(n1035), .Y(n1008) );
  BUFX2 U463 ( .A(n1034), .Y(n1012) );
  BUFX2 U464 ( .A(n1037), .Y(n1004) );
  BUFX2 U465 ( .A(n1037), .Y(n1003) );
  BUFX2 U466 ( .A(n1036), .Y(n1005) );
  BUFX2 U467 ( .A(n1032), .Y(n1017) );
  BUFX2 U468 ( .A(n1036), .Y(n1006) );
  BUFX2 U469 ( .A(n1034), .Y(n1011) );
  BUFX2 U470 ( .A(n1034), .Y(n1013) );
  BUFX2 U471 ( .A(n1033), .Y(n1014) );
  BUFX2 U472 ( .A(n1033), .Y(n1015) );
  BUFX2 U473 ( .A(n1035), .Y(n1009) );
  BUFX2 U474 ( .A(n1033), .Y(n1016) );
  BUFX2 U475 ( .A(n1035), .Y(n1010) );
  BUFX2 U476 ( .A(n1031), .Y(n1020) );
  BUFX2 U477 ( .A(n1031), .Y(n1021) );
  BUFX2 U478 ( .A(n1032), .Y(n1018) );
  BUFX2 U479 ( .A(n1032), .Y(n1019) );
  BUFX2 U480 ( .A(n1030), .Y(n1023) );
  BUFX2 U481 ( .A(n1030), .Y(n1024) );
  BUFX2 U482 ( .A(n1031), .Y(n1022) );
  BUFX2 U483 ( .A(n1029), .Y(n1027) );
  BUFX2 U484 ( .A(n1030), .Y(n1025) );
  BUFX2 U485 ( .A(n1029), .Y(n1026) );
  BUFX2 U486 ( .A(n916), .Y(n883) );
  BUFX2 U487 ( .A(n1857), .Y(n916) );
  BUFX2 U488 ( .A(n1029), .Y(n1028) );
  INVX2 U489 ( .A(n946), .Y(n936) );
  INVX2 U490 ( .A(n945), .Y(n934) );
  INVX2 U491 ( .A(n946), .Y(n933) );
  INVX2 U492 ( .A(n945), .Y(n932) );
  BUFX2 U493 ( .A(n948), .Y(n946) );
  BUFX2 U494 ( .A(n948), .Y(n945) );
  BUFX2 U495 ( .A(n880), .Y(n877) );
  BUFX2 U496 ( .A(n881), .Y(n876) );
  BUFX2 U497 ( .A(n881), .Y(n875) );
  BUFX2 U498 ( .A(n881), .Y(n874) );
  BUFX2 U499 ( .A(n880), .Y(n878) );
  BUFX2 U500 ( .A(n880), .Y(n879) );
  BUFX2 U501 ( .A(n1038), .Y(n1037) );
  BUFX2 U502 ( .A(n1038), .Y(n1036) );
  BUFX2 U503 ( .A(n1039), .Y(n1034) );
  BUFX2 U504 ( .A(n1039), .Y(n1033) );
  BUFX2 U505 ( .A(n1038), .Y(n1035) );
  BUFX2 U506 ( .A(n1039), .Y(n1032) );
  BUFX2 U507 ( .A(n1040), .Y(n1031) );
  BUFX2 U508 ( .A(n1040), .Y(n1030) );
  BUFX2 U509 ( .A(n1040), .Y(n1029) );
  BUFX2 U510 ( .A(n1000), .Y(n989) );
  BUFX2 U511 ( .A(n1000), .Y(n990) );
  BUFX2 U512 ( .A(n1000), .Y(n991) );
  BUFX2 U513 ( .A(n999), .Y(n992) );
  BUFX2 U514 ( .A(n999), .Y(n993) );
  BUFX2 U515 ( .A(n999), .Y(n994) );
  BUFX2 U516 ( .A(n998), .Y(n995) );
  BUFX2 U517 ( .A(n998), .Y(n996) );
  BUFX2 U518 ( .A(n1001), .Y(n987) );
  BUFX2 U519 ( .A(n1001), .Y(n988) );
  BUFX2 U520 ( .A(n337), .Y(n949) );
  BUFX2 U521 ( .A(n337), .Y(n950) );
  BUFX2 U522 ( .A(n998), .Y(n997) );
  BUFX2 U523 ( .A(n947), .Y(n951) );
  INVX2 U524 ( .A(n862), .Y(n855) );
  INVX2 U525 ( .A(n860), .Y(n856) );
  INVX2 U526 ( .A(n863), .Y(n854) );
  INVX2 U527 ( .A(n865), .Y(n853) );
  INVX2 U528 ( .A(n947), .Y(n935) );
  BUFX2 U529 ( .A(n948), .Y(n947) );
  BUFX2 U530 ( .A(n5081), .Y(n1000) );
  BUFX2 U531 ( .A(n5081), .Y(n999) );
  BUFX2 U532 ( .A(n5081), .Y(n998) );
  BUFX2 U533 ( .A(n5081), .Y(n1001) );
  BUFX2 U534 ( .A(n870), .Y(n864) );
  BUFX2 U535 ( .A(n870), .Y(n863) );
  BUFX2 U536 ( .A(n871), .Y(n862) );
  BUFX2 U537 ( .A(n871), .Y(n861) );
  BUFX2 U538 ( .A(n871), .Y(n860) );
  BUFX2 U539 ( .A(n872), .Y(n859) );
  BUFX2 U540 ( .A(n872), .Y(n858) );
  BUFX2 U541 ( .A(n872), .Y(n857) );
  BUFX2 U542 ( .A(n870), .Y(n865) );
  BUFX2 U543 ( .A(n869), .Y(n867) );
  BUFX2 U544 ( .A(n869), .Y(n866) );
  BUFX2 U545 ( .A(n1854), .Y(n881) );
  BUFX2 U546 ( .A(n1854), .Y(n880) );
  BUFX2 U547 ( .A(Inst_AEAD_u_cc_en_state), .Y(n1038) );
  BUFX2 U548 ( .A(Inst_AEAD_u_cc_en_state), .Y(n1039) );
  BUFX2 U549 ( .A(Inst_AEAD_u_cc_en_state), .Y(n1040) );
  BUFX2 U550 ( .A(n869), .Y(n868) );
  BUFX2 U551 ( .A(n982), .Y(n979) );
  BUFX2 U552 ( .A(n982), .Y(n980) );
  BUFX2 U553 ( .A(n882), .Y(n873) );
  BUFX2 U554 ( .A(n1854), .Y(n882) );
  BUFX2 U555 ( .A(n985), .Y(n970) );
  BUFX2 U556 ( .A(n985), .Y(n971) );
  BUFX2 U557 ( .A(n985), .Y(n972) );
  BUFX2 U558 ( .A(n984), .Y(n973) );
  BUFX2 U559 ( .A(n984), .Y(n974) );
  BUFX2 U560 ( .A(n984), .Y(n975) );
  BUFX2 U561 ( .A(n983), .Y(n976) );
  BUFX2 U562 ( .A(n983), .Y(n977) );
  BUFX2 U563 ( .A(n983), .Y(n978) );
  BUFX2 U564 ( .A(n337), .Y(n948) );
  BUFX2 U565 ( .A(n982), .Y(n981) );
  BUFX2 U566 ( .A(n1775), .Y(n869) );
  BUFX2 U567 ( .A(n1775), .Y(n871) );
  BUFX2 U568 ( .A(n1775), .Y(n872) );
  BUFX2 U569 ( .A(n1775), .Y(n870) );
  BUFX2 U570 ( .A(n5077), .Y(n985) );
  BUFX2 U571 ( .A(n5077), .Y(n984) );
  BUFX2 U572 ( .A(n5077), .Y(n983) );
  BUFX2 U573 ( .A(n5077), .Y(n982) );
  BUFX2 U574 ( .A(n986), .Y(n969) );
  BUFX2 U575 ( .A(n5077), .Y(n986) );
  INVX2 U576 ( .A(Inst_AEAD_u_input_sub_774_carry[5]), .Y(n1044) );
  INVX2 U577 ( .A(Inst_AEAD_u_input_sub_751_carry[14]), .Y(n1042) );
  XNOR2X1 U578 ( .A(Inst_AEAD_u_input_sgmt_len_15_), .B(
        Inst_AEAD_u_input_sub_751_carry[15]), .Y(Inst_AEAD_u_input_N143) );
  NAND2X2 U579 ( .A(n1041), .B(n1042), .Y(Inst_AEAD_u_input_sub_751_carry[15])
         );
  XNOR2X1 U580 ( .A(Inst_AEAD_u_input_sgmt_len_3_), .B(
        Inst_AEAD_u_input_sgmt_len_2_), .Y(Inst_AEAD_u_input_N131) );
  XNOR2X1 U581 ( .A(Inst_AEAD_u_input_sgmt_len_4_), .B(
        Inst_AEAD_u_input_sub_751_carry[4]), .Y(Inst_AEAD_u_input_N132) );
  XNOR2X1 U582 ( .A(Inst_AEAD_u_input_sgmt_len_5_), .B(
        Inst_AEAD_u_input_sub_751_carry[5]), .Y(Inst_AEAD_u_input_N133) );
  XNOR2X1 U583 ( .A(Inst_AEAD_u_input_sgmt_len_6_), .B(
        Inst_AEAD_u_input_sub_751_carry[6]), .Y(Inst_AEAD_u_input_N134) );
  XNOR2X1 U584 ( .A(Inst_AEAD_u_input_sgmt_len_7_), .B(
        Inst_AEAD_u_input_sub_751_carry[7]), .Y(Inst_AEAD_u_input_N135) );
  XNOR2X1 U585 ( .A(Inst_AEAD_u_input_sgmt_len_8_), .B(
        Inst_AEAD_u_input_sub_751_carry[8]), .Y(Inst_AEAD_u_input_N136) );
  XNOR2X1 U586 ( .A(Inst_AEAD_u_input_sgmt_len_9_), .B(
        Inst_AEAD_u_input_sub_751_carry[9]), .Y(Inst_AEAD_u_input_N137) );
  XNOR2X1 U587 ( .A(Inst_AEAD_u_input_sgmt_len_10_), .B(
        Inst_AEAD_u_input_sub_751_carry[10]), .Y(Inst_AEAD_u_input_N138) );
  XNOR2X1 U588 ( .A(Inst_AEAD_u_input_sgmt_len_11_), .B(
        Inst_AEAD_u_input_sub_751_carry[11]), .Y(Inst_AEAD_u_input_N139) );
  XNOR2X1 U589 ( .A(Inst_AEAD_u_input_sgmt_len_12_), .B(
        Inst_AEAD_u_input_sub_751_carry[12]), .Y(Inst_AEAD_u_input_N140) );
  XNOR2X1 U590 ( .A(Inst_AEAD_u_input_sgmt_len_13_), .B(
        Inst_AEAD_u_input_sub_751_carry[13]), .Y(Inst_AEAD_u_input_N141) );
  XNOR2X1 U591 ( .A(Inst_AEAD_u_input_sgmt_len_14_), .B(
        Inst_AEAD_u_input_sub_751_carry[14]), .Y(Inst_AEAD_u_input_N142) );
  XNOR2X1 U592 ( .A(Inst_AEAD_u_input_slen_6_), .B(
        Inst_AEAD_u_input_sub_774_carry[6]), .Y(Inst_AEAD_u_input_N220) );
  NAND2X2 U593 ( .A(n1043), .B(n1044), .Y(Inst_AEAD_u_input_sub_774_carry[6])
         );
  XNOR2X1 U594 ( .A(Inst_AEAD_u_input_slen_3_), .B(Inst_AEAD_u_input_slen_2_), 
        .Y(Inst_AEAD_u_input_N217) );
  XNOR2X1 U595 ( .A(Inst_AEAD_u_input_slen_4_), .B(
        Inst_AEAD_u_input_sub_774_carry[4]), .Y(Inst_AEAD_u_input_N218) );
  XNOR2X1 U596 ( .A(Inst_AEAD_u_input_slen_5_), .B(
        Inst_AEAD_u_input_sub_774_carry[5]), .Y(Inst_AEAD_u_input_N219) );
  OR2X2 U597 ( .A(Inst_AEAD_u_input_sgmt_len_4_), .B(
        Inst_AEAD_u_input_sub_751_carry[4]), .Y(
        Inst_AEAD_u_input_sub_751_carry[5]) );
  OR2X2 U598 ( .A(Inst_AEAD_u_input_sgmt_len_5_), .B(
        Inst_AEAD_u_input_sub_751_carry[5]), .Y(
        Inst_AEAD_u_input_sub_751_carry[6]) );
  OR2X2 U599 ( .A(Inst_AEAD_u_input_sgmt_len_6_), .B(
        Inst_AEAD_u_input_sub_751_carry[6]), .Y(
        Inst_AEAD_u_input_sub_751_carry[7]) );
  OR2X2 U600 ( .A(Inst_AEAD_u_input_sgmt_len_7_), .B(
        Inst_AEAD_u_input_sub_751_carry[7]), .Y(
        Inst_AEAD_u_input_sub_751_carry[8]) );
  OR2X2 U601 ( .A(Inst_AEAD_u_input_sgmt_len_8_), .B(
        Inst_AEAD_u_input_sub_751_carry[8]), .Y(
        Inst_AEAD_u_input_sub_751_carry[9]) );
  OR2X2 U602 ( .A(Inst_AEAD_u_input_sgmt_len_9_), .B(
        Inst_AEAD_u_input_sub_751_carry[9]), .Y(
        Inst_AEAD_u_input_sub_751_carry[10]) );
  OR2X2 U603 ( .A(Inst_AEAD_u_input_sgmt_len_10_), .B(
        Inst_AEAD_u_input_sub_751_carry[10]), .Y(
        Inst_AEAD_u_input_sub_751_carry[11]) );
  OR2X2 U604 ( .A(Inst_AEAD_u_input_sgmt_len_11_), .B(
        Inst_AEAD_u_input_sub_751_carry[11]), .Y(
        Inst_AEAD_u_input_sub_751_carry[12]) );
  OR2X2 U605 ( .A(Inst_AEAD_u_input_sgmt_len_12_), .B(
        Inst_AEAD_u_input_sub_751_carry[12]), .Y(
        Inst_AEAD_u_input_sub_751_carry[13]) );
  OR2X2 U606 ( .A(Inst_AEAD_u_input_slen_4_), .B(
        Inst_AEAD_u_input_sub_774_carry[4]), .Y(
        Inst_AEAD_u_input_sub_774_carry[5]) );
  OR2X2 U607 ( .A(Inst_AEAD_u_input_sgmt_len_13_), .B(
        Inst_AEAD_u_input_sub_751_carry[13]), .Y(
        Inst_AEAD_u_input_sub_751_carry[14]) );
  OR2X2 U608 ( .A(Inst_AEAD_u_input_sgmt_len_3_), .B(
        Inst_AEAD_u_input_sgmt_len_2_), .Y(Inst_AEAD_u_input_sub_751_carry[4])
         );
  OR2X2 U609 ( .A(Inst_AEAD_u_input_slen_3_), .B(Inst_AEAD_u_input_slen_2_), 
        .Y(Inst_AEAD_u_input_sub_774_carry[4]) );
  INVX2 U610 ( .A(Inst_AEAD_u_input_slen_5_), .Y(n1043) );
  INVX2 U611 ( .A(Inst_AEAD_u_input_sgmt_len_14_), .Y(n1041) );
  OAI31X1 U612 ( .A0(n1604), .A1(Inst_AEAD_u_input_ss_0_), .A2(n1605), .B0(
        Inst_AEAD_u_input_ss_1_), .Y(sdi_ready) );
  OAI2B1X1 U613 ( .A1N(n1606), .A0(Inst_AEAD_u_input_reg_sel_zero), .B0(n1607), 
        .Y(pdi_ready) );
  OAI21X1 U614 ( .A0(Inst_AEAD_u_input_n553), .A1(Inst_AEAD_u_input_n554), 
        .B0(Inst_AEAD_cmd_wr_ready), .Y(n1607) );
  AOI211X1 U615 ( .A0(n1608), .A1(n937), .B0(rst), .C0(n1609), .Y(n5072) );
  NOR2BX1 U616 ( .AN(Inst_AEAD_u_hdr_buffer_memory_1__18_), .B(n1611), .Y(
        n5075) );
  NOR2X1 U617 ( .A(n1612), .B(n1613), .Y(n5076) );
  OAI21X1 U618 ( .A0(n1614), .A1(n1615), .B0(n1616), .Y(n5078) );
  MXI2X1 U619 ( .A(Inst_AEAD_u_input_ploc_1_), .B(Inst_AEAD_bdi[15]), .S0(n471), .Y(n1616) );
  OAI21X1 U620 ( .A0(n1614), .A1(n1617), .B0(n1618), .Y(n5079) );
  MXI2X1 U621 ( .A(Inst_AEAD_u_input_ploc_0_), .B(Inst_AEAD_bdi[7]), .S0(n471), 
        .Y(n1618) );
  MX2X1 U622 ( .A(Inst_AEAD_u_input_vbytes_3_), .B(n1619), .S0(
        Inst_AEAD_u_input_n392), .Y(n5080) );
  CLKNAND2X2 U623 ( .A(n1620), .B(n1621), .Y(n5082) );
  MXI2X1 U624 ( .A(n1622), .B(n1623), .S0(Inst_AEAD_u_cc_u_cc_dp_rc_1_), .Y(
        n1620) );
  MXI2X1 U625 ( .A(n1624), .B(n1625), .S0(Inst_AEAD_u_cc_u_cc_dp_rc_0_), .Y(
        n5083) );
  OR2X1 U626 ( .A(n1626), .B(n1627), .Y(n1624) );
  MX2X1 U627 ( .A(n1628), .B(n1629), .S0(randd[0]), .Y(Inst_counter_n195) );
  AO22X1 U628 ( .A0(n1629), .A1(randd[1]), .B0(Inst_counter_N5), .B1(n1628), 
        .Y(Inst_counter_n194) );
  AO22X1 U629 ( .A0(n1629), .A1(randd[2]), .B0(Inst_counter_N6), .B1(n1628), 
        .Y(Inst_counter_n193) );
  AO22X1 U630 ( .A0(n1629), .A1(randd[3]), .B0(Inst_counter_N7), .B1(n1628), 
        .Y(Inst_counter_n192) );
  AO22X1 U631 ( .A0(n1629), .A1(randd[4]), .B0(Inst_counter_N8), .B1(n1628), 
        .Y(Inst_counter_n191) );
  AO22X1 U632 ( .A0(n1629), .A1(randd[5]), .B0(Inst_counter_N9), .B1(n1628), 
        .Y(Inst_counter_n190) );
  AO22X1 U633 ( .A0(n1629), .A1(randd[6]), .B0(Inst_counter_N10), .B1(n1628), 
        .Y(Inst_counter_n189) );
  AO22X1 U634 ( .A0(n1629), .A1(randd[7]), .B0(Inst_counter_N11), .B1(n1628), 
        .Y(Inst_counter_n188) );
  AO22X1 U635 ( .A0(n1629), .A1(randd[8]), .B0(Inst_counter_N12), .B1(n1628), 
        .Y(Inst_counter_n187) );
  AO22X1 U636 ( .A0(n1629), .A1(randd[9]), .B0(Inst_counter_N13), .B1(n1628), 
        .Y(Inst_counter_n186) );
  AO22X1 U637 ( .A0(n1629), .A1(randd[10]), .B0(Inst_counter_N14), .B1(n1628), 
        .Y(Inst_counter_n185) );
  AO22X1 U638 ( .A0(n1629), .A1(randd[11]), .B0(Inst_counter_N15), .B1(n1628), 
        .Y(Inst_counter_n184) );
  AO22X1 U639 ( .A0(n1629), .A1(randd[12]), .B0(Inst_counter_N16), .B1(n1628), 
        .Y(Inst_counter_n183) );
  AO22X1 U640 ( .A0(n1629), .A1(randd[13]), .B0(Inst_counter_N17), .B1(n1628), 
        .Y(Inst_counter_n182) );
  AO22X1 U641 ( .A0(n1629), .A1(randd[14]), .B0(Inst_counter_N18), .B1(n1628), 
        .Y(Inst_counter_n181) );
  AO22X1 U642 ( .A0(n1629), .A1(randd[15]), .B0(Inst_counter_N19), .B1(n1628), 
        .Y(Inst_counter_n180) );
  AO22X1 U643 ( .A0(n1629), .A1(randd[16]), .B0(Inst_counter_N20), .B1(n1628), 
        .Y(Inst_counter_n179) );
  AO22X1 U644 ( .A0(n1629), .A1(randd[17]), .B0(Inst_counter_N21), .B1(n1628), 
        .Y(Inst_counter_n178) );
  AO22X1 U645 ( .A0(n1629), .A1(randd[18]), .B0(Inst_counter_N22), .B1(n1628), 
        .Y(Inst_counter_n177) );
  AO22X1 U646 ( .A0(n1629), .A1(randd[19]), .B0(Inst_counter_N23), .B1(n1628), 
        .Y(Inst_counter_n176) );
  AO22X1 U647 ( .A0(n1629), .A1(randd[20]), .B0(Inst_counter_N24), .B1(n1628), 
        .Y(Inst_counter_n175) );
  AO22X1 U648 ( .A0(n1629), .A1(randd[21]), .B0(Inst_counter_N25), .B1(n1628), 
        .Y(Inst_counter_n174) );
  AO22X1 U649 ( .A0(n1629), .A1(randd[22]), .B0(Inst_counter_N26), .B1(n1628), 
        .Y(Inst_counter_n173) );
  AO22X1 U650 ( .A0(n1629), .A1(randd[23]), .B0(Inst_counter_N27), .B1(n1628), 
        .Y(Inst_counter_n172) );
  AO22X1 U651 ( .A0(n1629), .A1(randd[24]), .B0(Inst_counter_N28), .B1(n1628), 
        .Y(Inst_counter_n171) );
  AO22X1 U652 ( .A0(n1629), .A1(randd[25]), .B0(Inst_counter_N29), .B1(n1628), 
        .Y(Inst_counter_n170) );
  AO22X1 U653 ( .A0(n1629), .A1(randd[26]), .B0(Inst_counter_N30), .B1(n1628), 
        .Y(Inst_counter_n169) );
  AO22X1 U654 ( .A0(n1629), .A1(randd[27]), .B0(Inst_counter_N31), .B1(n1628), 
        .Y(Inst_counter_n168) );
  AO22X1 U655 ( .A0(n1629), .A1(randd[28]), .B0(Inst_counter_N32), .B1(n1628), 
        .Y(Inst_counter_n167) );
  AO22X1 U656 ( .A0(n1629), .A1(randd[29]), .B0(Inst_counter_N33), .B1(n1628), 
        .Y(Inst_counter_n166) );
  AO22X1 U657 ( .A0(n1629), .A1(randd[30]), .B0(Inst_counter_N34), .B1(n1628), 
        .Y(Inst_counter_n165) );
  AO22X1 U658 ( .A0(n1629), .A1(randd[31]), .B0(Inst_counter_N35), .B1(n1628), 
        .Y(Inst_counter_n164) );
  AO22X1 U659 ( .A0(n1629), .A1(randd[32]), .B0(Inst_counter_N36), .B1(n1628), 
        .Y(Inst_counter_n163) );
  AO22X1 U660 ( .A0(n1629), .A1(randd[33]), .B0(Inst_counter_N37), .B1(n1628), 
        .Y(Inst_counter_n162) );
  AO22X1 U661 ( .A0(n1629), .A1(randd[34]), .B0(Inst_counter_N38), .B1(n1628), 
        .Y(Inst_counter_n161) );
  AO22X1 U662 ( .A0(n1629), .A1(randd[35]), .B0(Inst_counter_N39), .B1(n1628), 
        .Y(Inst_counter_n160) );
  AO22X1 U663 ( .A0(n1629), .A1(randd[36]), .B0(Inst_counter_N40), .B1(n1628), 
        .Y(Inst_counter_n159) );
  AO22X1 U664 ( .A0(n1629), .A1(randd[37]), .B0(Inst_counter_N41), .B1(n1628), 
        .Y(Inst_counter_n158) );
  AO22X1 U665 ( .A0(n1629), .A1(randd[38]), .B0(Inst_counter_N42), .B1(n1628), 
        .Y(Inst_counter_n157) );
  AO22X1 U666 ( .A0(n1629), .A1(randd[39]), .B0(Inst_counter_N43), .B1(n1628), 
        .Y(Inst_counter_n156) );
  AO22X1 U667 ( .A0(n1629), .A1(randd[40]), .B0(Inst_counter_N44), .B1(n1628), 
        .Y(Inst_counter_n155) );
  AO22X1 U668 ( .A0(n1629), .A1(randd[41]), .B0(Inst_counter_N45), .B1(n1628), 
        .Y(Inst_counter_n154) );
  AO22X1 U669 ( .A0(n1629), .A1(randd[42]), .B0(Inst_counter_N46), .B1(n1628), 
        .Y(Inst_counter_n153) );
  AO22X1 U670 ( .A0(n1629), .A1(randd[43]), .B0(Inst_counter_N47), .B1(n1628), 
        .Y(Inst_counter_n152) );
  AO22X1 U671 ( .A0(n1629), .A1(randd[44]), .B0(Inst_counter_N48), .B1(n1628), 
        .Y(Inst_counter_n151) );
  AO22X1 U672 ( .A0(n1629), .A1(randd[45]), .B0(Inst_counter_N49), .B1(n1628), 
        .Y(Inst_counter_n150) );
  AO22X1 U673 ( .A0(n1629), .A1(randd[46]), .B0(Inst_counter_N50), .B1(n1628), 
        .Y(Inst_counter_n149) );
  AO22X1 U674 ( .A0(n1629), .A1(randd[47]), .B0(Inst_counter_N51), .B1(n1628), 
        .Y(Inst_counter_n148) );
  AO22X1 U675 ( .A0(n1629), .A1(randd[48]), .B0(Inst_counter_N52), .B1(n1628), 
        .Y(Inst_counter_n147) );
  AO22X1 U676 ( .A0(n1629), .A1(randd[49]), .B0(Inst_counter_N53), .B1(n1628), 
        .Y(Inst_counter_n146) );
  AO22X1 U677 ( .A0(n1629), .A1(randd[50]), .B0(Inst_counter_N54), .B1(n1628), 
        .Y(Inst_counter_n145) );
  AO22X1 U678 ( .A0(n1629), .A1(randd[51]), .B0(Inst_counter_N55), .B1(n1628), 
        .Y(Inst_counter_n144) );
  AO22X1 U679 ( .A0(n1629), .A1(randd[52]), .B0(Inst_counter_N56), .B1(n1628), 
        .Y(Inst_counter_n143) );
  AO22X1 U680 ( .A0(n1629), .A1(randd[53]), .B0(Inst_counter_N57), .B1(n1628), 
        .Y(Inst_counter_n142) );
  AO22X1 U681 ( .A0(n1629), .A1(randd[54]), .B0(Inst_counter_N58), .B1(n1628), 
        .Y(Inst_counter_n141) );
  AO22X1 U682 ( .A0(n1629), .A1(randd[55]), .B0(Inst_counter_N59), .B1(n1628), 
        .Y(Inst_counter_n140) );
  AO22X1 U683 ( .A0(n1629), .A1(randd[56]), .B0(Inst_counter_N60), .B1(n1628), 
        .Y(Inst_counter_n139) );
  AO22X1 U684 ( .A0(n1629), .A1(randd[57]), .B0(Inst_counter_N61), .B1(n1628), 
        .Y(Inst_counter_n138) );
  AO22X1 U685 ( .A0(n1629), .A1(randd[58]), .B0(Inst_counter_N62), .B1(n1628), 
        .Y(Inst_counter_n137) );
  AO22X1 U686 ( .A0(n1629), .A1(randd[59]), .B0(Inst_counter_N63), .B1(n1628), 
        .Y(Inst_counter_n136) );
  AO22X1 U687 ( .A0(n1629), .A1(randd[60]), .B0(Inst_counter_N64), .B1(n1628), 
        .Y(Inst_counter_n135) );
  AO22X1 U688 ( .A0(n1629), .A1(randd[61]), .B0(Inst_counter_N65), .B1(n1628), 
        .Y(Inst_counter_n134) );
  AO22X1 U689 ( .A0(n1629), .A1(randd[62]), .B0(Inst_counter_N66), .B1(n1628), 
        .Y(Inst_counter_n133) );
  MXI2X1 U690 ( .A(n1630), .B(n1631), .S0(randd[63]), .Y(Inst_counter_n132) );
  AOI2B1X1 U691 ( .A1N(Inst_counter_add_3021_carry[63]), .A0(n1628), .B0(n1629), .Y(n1631) );
  CLKNAND2X2 U692 ( .A(Inst_counter_add_3021_carry[63]), .B(n1628), .Y(n1630)
         );
  MX2X1 U693 ( .A(IDtReg[48]), .B(IDt[48]), .S0(ld_rec), .Y(Inst_RegIDt_n99)
         );
  MX2X1 U694 ( .A(IDtReg[47]), .B(IDt[47]), .S0(ld_rec), .Y(Inst_RegIDt_n97)
         );
  MX2X1 U695 ( .A(IDtReg[46]), .B(IDt[46]), .S0(ld_rec), .Y(Inst_RegIDt_n95)
         );
  MX2X1 U696 ( .A(IDtReg[45]), .B(IDt[45]), .S0(ld_rec), .Y(Inst_RegIDt_n93)
         );
  MX2X1 U697 ( .A(IDtReg[44]), .B(IDt[44]), .S0(ld_rec), .Y(Inst_RegIDt_n91)
         );
  MX2X1 U698 ( .A(IDtReg[3]), .B(IDt[3]), .S0(ld_rec), .Y(Inst_RegIDt_n9) );
  MX2X1 U699 ( .A(IDtReg[43]), .B(IDt[43]), .S0(ld_rec), .Y(Inst_RegIDt_n89)
         );
  MX2X1 U700 ( .A(IDtReg[42]), .B(IDt[42]), .S0(ld_rec), .Y(Inst_RegIDt_n87)
         );
  MX2X1 U701 ( .A(IDtReg[41]), .B(IDt[41]), .S0(ld_rec), .Y(Inst_RegIDt_n85)
         );
  MX2X1 U702 ( .A(IDtReg[40]), .B(IDt[40]), .S0(ld_rec), .Y(Inst_RegIDt_n83)
         );
  MX2X1 U703 ( .A(IDtReg[39]), .B(IDt[39]), .S0(ld_rec), .Y(Inst_RegIDt_n81)
         );
  MX2X1 U704 ( .A(IDtReg[38]), .B(IDt[38]), .S0(ld_rec), .Y(Inst_RegIDt_n79)
         );
  MX2X1 U705 ( .A(IDtReg[37]), .B(IDt[37]), .S0(ld_rec), .Y(Inst_RegIDt_n77)
         );
  MX2X1 U706 ( .A(IDtReg[36]), .B(IDt[36]), .S0(ld_rec), .Y(Inst_RegIDt_n75)
         );
  MX2X1 U707 ( .A(IDtReg[35]), .B(IDt[35]), .S0(ld_rec), .Y(Inst_RegIDt_n73)
         );
  MX2X1 U708 ( .A(IDtReg[34]), .B(IDt[34]), .S0(ld_rec), .Y(Inst_RegIDt_n71)
         );
  MX2X1 U709 ( .A(IDtReg[2]), .B(IDt[2]), .S0(ld_rec), .Y(Inst_RegIDt_n7) );
  MX2X1 U710 ( .A(IDtReg[33]), .B(IDt[33]), .S0(ld_rec), .Y(Inst_RegIDt_n69)
         );
  MX2X1 U711 ( .A(IDtReg[32]), .B(IDt[32]), .S0(ld_rec), .Y(Inst_RegIDt_n67)
         );
  MX2X1 U712 ( .A(IDtReg[31]), .B(IDt[31]), .S0(ld_rec), .Y(Inst_RegIDt_n65)
         );
  MX2X1 U713 ( .A(IDtReg[30]), .B(IDt[30]), .S0(ld_rec), .Y(Inst_RegIDt_n63)
         );
  MX2X1 U714 ( .A(IDtReg[29]), .B(IDt[29]), .S0(ld_rec), .Y(Inst_RegIDt_n61)
         );
  MX2X1 U715 ( .A(IDtReg[28]), .B(IDt[28]), .S0(ld_rec), .Y(Inst_RegIDt_n59)
         );
  MX2X1 U716 ( .A(IDtReg[27]), .B(IDt[27]), .S0(ld_rec), .Y(Inst_RegIDt_n57)
         );
  MX2X1 U717 ( .A(IDtReg[26]), .B(IDt[26]), .S0(ld_rec), .Y(Inst_RegIDt_n55)
         );
  MX2X1 U718 ( .A(IDtReg[25]), .B(IDt[25]), .S0(ld_rec), .Y(Inst_RegIDt_n53)
         );
  MX2X1 U719 ( .A(IDtReg[24]), .B(IDt[24]), .S0(ld_rec), .Y(Inst_RegIDt_n51)
         );
  MX2X1 U720 ( .A(IDtReg[1]), .B(IDt[1]), .S0(ld_rec), .Y(Inst_RegIDt_n5) );
  MX2X1 U721 ( .A(IDtReg[23]), .B(IDt[23]), .S0(ld_rec), .Y(Inst_RegIDt_n49)
         );
  MX2X1 U722 ( .A(IDtReg[22]), .B(IDt[22]), .S0(ld_rec), .Y(Inst_RegIDt_n47)
         );
  MX2X1 U723 ( .A(IDtReg[21]), .B(IDt[21]), .S0(ld_rec), .Y(Inst_RegIDt_n45)
         );
  MX2X1 U724 ( .A(IDtReg[20]), .B(IDt[20]), .S0(ld_rec), .Y(Inst_RegIDt_n43)
         );
  MX2X1 U725 ( .A(IDtReg[19]), .B(IDt[19]), .S0(ld_rec), .Y(Inst_RegIDt_n41)
         );
  MX2X1 U726 ( .A(IDtReg[18]), .B(IDt[18]), .S0(ld_rec), .Y(Inst_RegIDt_n39)
         );
  MX2X1 U727 ( .A(IDtReg[17]), .B(IDt[17]), .S0(ld_rec), .Y(Inst_RegIDt_n37)
         );
  MX2X1 U728 ( .A(IDtReg[16]), .B(IDt[16]), .S0(ld_rec), .Y(Inst_RegIDt_n35)
         );
  MX2X1 U729 ( .A(IDtReg[15]), .B(IDt[15]), .S0(ld_rec), .Y(Inst_RegIDt_n33)
         );
  MX2X1 U730 ( .A(IDtReg[14]), .B(IDt[14]), .S0(ld_rec), .Y(Inst_RegIDt_n31)
         );
  MX2X1 U731 ( .A(IDtReg[0]), .B(IDt[0]), .S0(ld_rec), .Y(Inst_RegIDt_n3) );
  MX2X1 U732 ( .A(IDtReg[13]), .B(IDt[13]), .S0(ld_rec), .Y(Inst_RegIDt_n29)
         );
  MX2X1 U733 ( .A(IDtReg[12]), .B(IDt[12]), .S0(ld_rec), .Y(Inst_RegIDt_n27)
         );
  MX2X1 U734 ( .A(IDtReg[11]), .B(IDt[11]), .S0(ld_rec), .Y(Inst_RegIDt_n25)
         );
  MX2X1 U735 ( .A(IDtReg[10]), .B(IDt[10]), .S0(ld_rec), .Y(Inst_RegIDt_n23)
         );
  MX2X1 U736 ( .A(IDtReg[9]), .B(IDt[9]), .S0(ld_rec), .Y(Inst_RegIDt_n21) );
  MX2X1 U737 ( .A(IDtReg[8]), .B(IDt[8]), .S0(ld_rec), .Y(Inst_RegIDt_n19) );
  MX2X1 U738 ( .A(IDtReg[7]), .B(IDt[7]), .S0(ld_rec), .Y(Inst_RegIDt_n17) );
  MX2X1 U739 ( .A(IDtReg[6]), .B(IDt[6]), .S0(ld_rec), .Y(Inst_RegIDt_n15) );
  MX2X1 U740 ( .A(IDtReg[63]), .B(IDt[63]), .S0(ld_rec), .Y(Inst_RegIDt_n130)
         );
  MX2X1 U741 ( .A(IDtReg[5]), .B(IDt[5]), .S0(ld_rec), .Y(Inst_RegIDt_n13) );
  MX2X1 U742 ( .A(IDtReg[62]), .B(IDt[62]), .S0(ld_rec), .Y(Inst_RegIDt_n127)
         );
  MX2X1 U743 ( .A(IDtReg[61]), .B(IDt[61]), .S0(ld_rec), .Y(Inst_RegIDt_n125)
         );
  MX2X1 U744 ( .A(IDtReg[60]), .B(IDt[60]), .S0(ld_rec), .Y(Inst_RegIDt_n123)
         );
  MX2X1 U745 ( .A(IDtReg[59]), .B(IDt[59]), .S0(ld_rec), .Y(Inst_RegIDt_n121)
         );
  MX2X1 U746 ( .A(IDtReg[58]), .B(IDt[58]), .S0(ld_rec), .Y(Inst_RegIDt_n119)
         );
  MX2X1 U747 ( .A(IDtReg[57]), .B(IDt[57]), .S0(ld_rec), .Y(Inst_RegIDt_n117)
         );
  MX2X1 U748 ( .A(IDtReg[56]), .B(IDt[56]), .S0(ld_rec), .Y(Inst_RegIDt_n115)
         );
  MX2X1 U749 ( .A(IDtReg[55]), .B(IDt[55]), .S0(ld_rec), .Y(Inst_RegIDt_n113)
         );
  MX2X1 U750 ( .A(IDtReg[54]), .B(IDt[54]), .S0(ld_rec), .Y(Inst_RegIDt_n111)
         );
  MX2X1 U751 ( .A(IDtReg[4]), .B(IDt[4]), .S0(ld_rec), .Y(Inst_RegIDt_n11) );
  MX2X1 U752 ( .A(IDtReg[53]), .B(IDt[53]), .S0(ld_rec), .Y(Inst_RegIDt_n109)
         );
  MX2X1 U753 ( .A(IDtReg[52]), .B(IDt[52]), .S0(ld_rec), .Y(Inst_RegIDt_n107)
         );
  MX2X1 U754 ( .A(IDtReg[51]), .B(IDt[51]), .S0(ld_rec), .Y(Inst_RegIDt_n105)
         );
  MX2X1 U755 ( .A(IDtReg[50]), .B(IDt[50]), .S0(ld_rec), .Y(Inst_RegIDt_n103)
         );
  MX2X1 U756 ( .A(IDtReg[49]), .B(IDt[49]), .S0(ld_rec), .Y(Inst_RegIDt_n101)
         );
  MX2X1 U757 ( .A(IDstReg[48]), .B(IDst[48]), .S0(ld_rec), .Y(n5184) );
  MX2X1 U758 ( .A(IDstReg[47]), .B(IDst[47]), .S0(ld_rec), .Y(n5182) );
  MX2X1 U759 ( .A(IDstReg[46]), .B(IDst[46]), .S0(ld_rec), .Y(n5180) );
  MX2X1 U760 ( .A(IDstReg[45]), .B(IDst[45]), .S0(ld_rec), .Y(n5178) );
  MX2X1 U761 ( .A(IDstReg[44]), .B(IDst[44]), .S0(ld_rec), .Y(n5176) );
  MX2X1 U762 ( .A(IDstReg[3]), .B(IDst[3]), .S0(ld_rec), .Y(n5094) );
  MX2X1 U763 ( .A(IDstReg[43]), .B(IDst[43]), .S0(ld_rec), .Y(n5174) );
  MX2X1 U764 ( .A(IDstReg[42]), .B(IDst[42]), .S0(ld_rec), .Y(n5172) );
  MX2X1 U765 ( .A(IDstReg[41]), .B(IDst[41]), .S0(ld_rec), .Y(n5170) );
  MX2X1 U766 ( .A(IDstReg[40]), .B(IDst[40]), .S0(ld_rec), .Y(n5168) );
  MX2X1 U767 ( .A(IDstReg[39]), .B(IDst[39]), .S0(ld_rec), .Y(n5166) );
  MX2X1 U768 ( .A(IDstReg[38]), .B(IDst[38]), .S0(ld_rec), .Y(n5164) );
  MX2X1 U769 ( .A(IDstReg[37]), .B(IDst[37]), .S0(ld_rec), .Y(n5162) );
  MX2X1 U770 ( .A(IDstReg[36]), .B(IDst[36]), .S0(ld_rec), .Y(n5160) );
  MX2X1 U771 ( .A(IDstReg[35]), .B(IDst[35]), .S0(ld_rec), .Y(n5158) );
  MX2X1 U772 ( .A(IDstReg[34]), .B(IDst[34]), .S0(ld_rec), .Y(n5156) );
  MX2X1 U773 ( .A(IDstReg[2]), .B(IDst[2]), .S0(ld_rec), .Y(n5092) );
  MX2X1 U774 ( .A(IDstReg[33]), .B(IDst[33]), .S0(ld_rec), .Y(n5154) );
  MX2X1 U775 ( .A(IDstReg[32]), .B(IDst[32]), .S0(ld_rec), .Y(n5152) );
  MX2X1 U776 ( .A(IDstReg[31]), .B(IDst[31]), .S0(ld_rec), .Y(n5150) );
  MX2X1 U777 ( .A(IDstReg[30]), .B(IDst[30]), .S0(ld_rec), .Y(n5148) );
  MX2X1 U778 ( .A(IDstReg[29]), .B(IDst[29]), .S0(ld_rec), .Y(n5146) );
  MX2X1 U779 ( .A(IDstReg[28]), .B(IDst[28]), .S0(ld_rec), .Y(n5144) );
  MX2X1 U780 ( .A(IDstReg[27]), .B(IDst[27]), .S0(ld_rec), .Y(n5142) );
  MX2X1 U781 ( .A(IDstReg[26]), .B(IDst[26]), .S0(ld_rec), .Y(n5140) );
  MX2X1 U782 ( .A(IDstReg[25]), .B(IDst[25]), .S0(ld_rec), .Y(n5138) );
  MX2X1 U783 ( .A(IDstReg[24]), .B(IDst[24]), .S0(ld_rec), .Y(n5136) );
  MX2X1 U784 ( .A(IDstReg[1]), .B(IDst[1]), .S0(ld_rec), .Y(n5090) );
  MX2X1 U785 ( .A(IDstReg[23]), .B(IDst[23]), .S0(ld_rec), .Y(n5134) );
  MX2X1 U786 ( .A(IDstReg[22]), .B(IDst[22]), .S0(ld_rec), .Y(n5132) );
  MX2X1 U787 ( .A(IDstReg[21]), .B(IDst[21]), .S0(ld_rec), .Y(n5130) );
  MX2X1 U788 ( .A(IDstReg[20]), .B(IDst[20]), .S0(ld_rec), .Y(n5128) );
  MX2X1 U789 ( .A(IDstReg[19]), .B(IDst[19]), .S0(ld_rec), .Y(n5126) );
  MX2X1 U790 ( .A(IDstReg[18]), .B(IDst[18]), .S0(ld_rec), .Y(n5124) );
  MX2X1 U791 ( .A(IDstReg[17]), .B(IDst[17]), .S0(ld_rec), .Y(n5122) );
  MX2X1 U792 ( .A(IDstReg[16]), .B(IDst[16]), .S0(ld_rec), .Y(n5120) );
  MX2X1 U793 ( .A(IDstReg[15]), .B(IDst[15]), .S0(ld_rec), .Y(n5118) );
  MX2X1 U794 ( .A(IDstReg[14]), .B(IDst[14]), .S0(ld_rec), .Y(n5116) );
  MX2X1 U795 ( .A(IDstReg[0]), .B(IDst[0]), .S0(ld_rec), .Y(n5088) );
  MX2X1 U796 ( .A(IDstReg[13]), .B(IDst[13]), .S0(ld_rec), .Y(n5114) );
  MX2X1 U797 ( .A(IDstReg[12]), .B(IDst[12]), .S0(ld_rec), .Y(n5112) );
  MX2X1 U798 ( .A(IDstReg[11]), .B(IDst[11]), .S0(ld_rec), .Y(n5110) );
  MX2X1 U799 ( .A(IDstReg[10]), .B(IDst[10]), .S0(ld_rec), .Y(n5108) );
  MX2X1 U800 ( .A(IDstReg[9]), .B(IDst[9]), .S0(ld_rec), .Y(n5106) );
  MX2X1 U801 ( .A(IDstReg[8]), .B(IDst[8]), .S0(ld_rec), .Y(n5104) );
  MX2X1 U802 ( .A(IDstReg[7]), .B(IDst[7]), .S0(ld_rec), .Y(n5102) );
  MX2X1 U803 ( .A(IDstReg[6]), .B(IDst[6]), .S0(ld_rec), .Y(n5100) );
  MX2X1 U804 ( .A(IDstReg[63]), .B(IDst[63]), .S0(ld_rec), .Y(n5214) );
  MX2X1 U805 ( .A(IDstReg[5]), .B(IDst[5]), .S0(ld_rec), .Y(n5098) );
  MX2X1 U806 ( .A(IDstReg[62]), .B(IDst[62]), .S0(ld_rec), .Y(n5212) );
  MX2X1 U807 ( .A(IDstReg[61]), .B(IDst[61]), .S0(ld_rec), .Y(n5210) );
  MX2X1 U808 ( .A(IDstReg[60]), .B(IDst[60]), .S0(ld_rec), .Y(n5208) );
  MX2X1 U809 ( .A(IDstReg[59]), .B(IDst[59]), .S0(ld_rec), .Y(n5206) );
  MX2X1 U810 ( .A(IDstReg[58]), .B(IDst[58]), .S0(ld_rec), .Y(n5204) );
  MX2X1 U811 ( .A(IDstReg[57]), .B(IDst[57]), .S0(ld_rec), .Y(n5202) );
  MX2X1 U812 ( .A(IDstReg[56]), .B(IDst[56]), .S0(ld_rec), .Y(n5200) );
  MX2X1 U813 ( .A(IDstReg[55]), .B(IDst[55]), .S0(ld_rec), .Y(n5198) );
  MX2X1 U814 ( .A(IDstReg[54]), .B(IDst[54]), .S0(ld_rec), .Y(n5196) );
  MX2X1 U815 ( .A(IDstReg[4]), .B(IDst[4]), .S0(ld_rec), .Y(n5096) );
  MX2X1 U816 ( .A(IDstReg[53]), .B(IDst[53]), .S0(ld_rec), .Y(n5194) );
  MX2X1 U817 ( .A(IDstReg[52]), .B(IDst[52]), .S0(ld_rec), .Y(n5192) );
  MX2X1 U818 ( .A(IDstReg[51]), .B(IDst[51]), .S0(ld_rec), .Y(n5190) );
  MX2X1 U819 ( .A(IDstReg[50]), .B(IDst[50]), .S0(ld_rec), .Y(n5188) );
  MX2X1 U820 ( .A(IDstReg[49]), .B(IDst[49]), .S0(ld_rec), .Y(n5186) );
  OAI2B2X1 U821 ( .A1N(Inst_AEAD_key[0]), .A0(n1632), .B0(
        Inst_AEAD_u_input_n362), .B1(n1633), .Y(Inst_AEAD_u_input_n552) );
  OAI2B1X1 U822 ( .A1N(Inst_AEAD_key[6]), .A0(n1632), .B0(n1634), .Y(
        Inst_AEAD_u_input_n551) );
  AOI22XL U823 ( .A0(Inst_AEAD_u_input_N220), .A1(n1635), .B0(
        Inst_AEAD_u_input_slen_6_), .B1(n1636), .Y(n1634) );
  OAI32XL U824 ( .A0(n1632), .A1(rst), .A2(n1637), .B0(n1638), .B1(n1639), .Y(
        Inst_AEAD_u_input_n550) );
  AOI21X1 U825 ( .A0(n981), .A1(n1640), .B0(n1637), .Y(n1638) );
  NAND4X1 U826 ( .A(Inst_AEAD_u_input_n362), .B(n466), .C(
        Inst_AEAD_u_input_slen_2_), .D(n1641), .Y(n1640) );
  NOR4X1 U827 ( .A(Inst_AEAD_u_input_slen_6_), .B(Inst_AEAD_u_input_slen_5_), 
        .C(Inst_AEAD_u_input_slen_4_), .D(Inst_AEAD_u_input_slen_3_), .Y(n1641) );
  MX2X1 U828 ( .A(n1642), .B(n1637), .S0(Inst_AEAD_u_input_ss_0_), .Y(
        Inst_AEAD_u_input_n549) );
  NOR4BX1 U829 ( .AN(n1643), .B(Inst_AEAD_key[29]), .C(Inst_AEAD_key[31]), .D(
        Inst_AEAD_key[28]), .Y(n1642) );
  NOR4BX1 U830 ( .AN(Inst_AEAD_key[30]), .B(rst), .C(Inst_AEAD_u_input_ss_1_), 
        .D(n1637), .Y(n1643) );
  AND2X1 U831 ( .A(n1644), .B(n981), .Y(n1637) );
  MXI2X1 U832 ( .A(n1645), .B(sdi_valid), .S0(n1639), .Y(n1644) );
  AOI2BB1X1 U833 ( .A0N(Inst_AEAD_u_input_ss_0_), .A1N(sdi_valid), .B0(n1605), 
        .Y(n1645) );
  OAI2B2X1 U834 ( .A1N(Inst_AEAD_key[1]), .A0(n1632), .B0(n1633), .B1(n466), 
        .Y(Inst_AEAD_u_input_n548) );
  NOR2X1 U835 ( .A(n1636), .B(n1635), .Y(n1633) );
  OAI2B1X1 U836 ( .A1N(Inst_AEAD_key[2]), .A0(n1632), .B0(n1646), .Y(
        Inst_AEAD_u_input_n547) );
  MXI2X1 U837 ( .A(n1635), .B(n1636), .S0(Inst_AEAD_u_input_slen_2_), .Y(n1646) );
  OAI2B1X1 U838 ( .A1N(Inst_AEAD_key[3]), .A0(n1632), .B0(n1647), .Y(
        Inst_AEAD_u_input_n546) );
  AOI22XL U839 ( .A0(Inst_AEAD_u_input_N217), .A1(n1635), .B0(
        Inst_AEAD_u_input_slen_3_), .B1(n1636), .Y(n1647) );
  OAI2B1X1 U840 ( .A1N(Inst_AEAD_key[4]), .A0(n1632), .B0(n1648), .Y(
        Inst_AEAD_u_input_n545) );
  AOI22XL U841 ( .A0(Inst_AEAD_u_input_N218), .A1(n1635), .B0(
        Inst_AEAD_u_input_slen_4_), .B1(n1636), .Y(n1648) );
  OAI2B1X1 U842 ( .A1N(Inst_AEAD_key[5]), .A0(n1632), .B0(n1649), .Y(
        Inst_AEAD_u_input_n544) );
  AOI22XL U843 ( .A0(Inst_AEAD_u_input_N219), .A1(n1635), .B0(
        Inst_AEAD_u_input_slen_5_), .B1(n1636), .Y(n1649) );
  NOR2BX1 U844 ( .AN(n1632), .B(n1636), .Y(n1635) );
  OA21X1 U845 ( .A0(n1605), .A1(n1650), .B0(n1632), .Y(n1636) );
  OAI21X1 U846 ( .A0(Inst_AEAD_u_input_ss_0_), .A1(sdi_valid), .B0(
        Inst_AEAD_u_input_ss_1_), .Y(n1650) );
  CLKNAND2X2 U847 ( .A(Inst_AEAD_u_input_ss_0_), .B(n1639), .Y(n1632) );
  NOR3X1 U848 ( .A(n1651), .B(Inst_AEAD_u_input_n553), .C(n1652), .Y(
        Inst_AEAD_u_input_n543) );
  XNOR2X1 U849 ( .A(n472), .B(Inst_AEAD_u_input_ctr_0_), .Y(n1651) );
  NOR3BX1 U850 ( .AN(n1653), .B(n1654), .C(Inst_AEAD_u_input_n554), .Y(
        Inst_AEAD_u_input_n542) );
  OAI22X1 U851 ( .A0(rst), .A1(n1655), .B0(n1656), .B1(n1657), .Y(
        Inst_AEAD_u_input_n541) );
  OAI21X1 U852 ( .A0(n5086), .A1(n1615), .B0(n1658), .Y(Inst_AEAD_u_input_n540) );
  AOI22XL U853 ( .A0(Inst_AEAD_u_input_N143), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_15_), .B1(n1660), .Y(n1658) );
  OAI22X1 U854 ( .A0(n5086), .A1(n1661), .B0(n1662), .B1(n1663), .Y(
        Inst_AEAD_u_input_n539) );
  OAI22X1 U855 ( .A0(n5086), .A1(n1664), .B0(n1662), .B1(n1665), .Y(
        Inst_AEAD_u_input_n538) );
  NOR2X1 U856 ( .A(n1660), .B(n1659), .Y(n1662) );
  OAI21X1 U857 ( .A0(n5086), .A1(n1666), .B0(n1667), .Y(Inst_AEAD_u_input_n537) );
  MXI2X1 U858 ( .A(n1659), .B(n1660), .S0(Inst_AEAD_u_input_sgmt_len_2_), .Y(
        n1667) );
  OAI21X1 U859 ( .A0(n5086), .A1(n1668), .B0(n1669), .Y(Inst_AEAD_u_input_n536) );
  AOI22XL U860 ( .A0(Inst_AEAD_u_input_N131), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_3_), .B1(n1660), .Y(n1669) );
  OAI21X1 U861 ( .A0(n5086), .A1(n1670), .B0(n1671), .Y(Inst_AEAD_u_input_n535) );
  AOI22XL U862 ( .A0(Inst_AEAD_u_input_N132), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_4_), .B1(n1660), .Y(n1671) );
  OAI21X1 U863 ( .A0(n5086), .A1(n1672), .B0(n1673), .Y(Inst_AEAD_u_input_n534) );
  AOI22XL U864 ( .A0(Inst_AEAD_u_input_N133), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_5_), .B1(n1660), .Y(n1673) );
  OAI21X1 U865 ( .A0(n5086), .A1(n1674), .B0(n1675), .Y(Inst_AEAD_u_input_n533) );
  AOI22XL U866 ( .A0(Inst_AEAD_u_input_N134), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_6_), .B1(n1660), .Y(n1675) );
  OAI21X1 U867 ( .A0(n5086), .A1(n1617), .B0(n1676), .Y(Inst_AEAD_u_input_n532) );
  AOI22XL U868 ( .A0(Inst_AEAD_u_input_N135), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_7_), .B1(n1660), .Y(n1676) );
  OAI21X1 U869 ( .A0(n5086), .A1(n1677), .B0(n1678), .Y(Inst_AEAD_u_input_n531) );
  AOI22XL U870 ( .A0(Inst_AEAD_u_input_N136), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_8_), .B1(n1660), .Y(n1678) );
  OAI21X1 U871 ( .A0(n5086), .A1(n1679), .B0(n1680), .Y(Inst_AEAD_u_input_n530) );
  AOI22XL U872 ( .A0(Inst_AEAD_u_input_N137), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_9_), .B1(n1660), .Y(n1680) );
  OAI21X1 U873 ( .A0(n5086), .A1(n1681), .B0(n1682), .Y(Inst_AEAD_u_input_n529) );
  AOI22XL U874 ( .A0(Inst_AEAD_u_input_N138), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_10_), .B1(n1660), .Y(n1682) );
  OAI21X1 U875 ( .A0(n5086), .A1(n1683), .B0(n1684), .Y(Inst_AEAD_u_input_n528) );
  AOI22XL U876 ( .A0(Inst_AEAD_u_input_N139), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_11_), .B1(n1660), .Y(n1684) );
  OAI21X1 U877 ( .A0(n5086), .A1(n1685), .B0(n1686), .Y(Inst_AEAD_u_input_n527) );
  AOI22XL U878 ( .A0(Inst_AEAD_u_input_N140), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_12_), .B1(n1660), .Y(n1686) );
  OAI21X1 U879 ( .A0(n5086), .A1(n1687), .B0(n1688), .Y(Inst_AEAD_u_input_n526) );
  AOI22XL U880 ( .A0(Inst_AEAD_u_input_N141), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_13_), .B1(n1660), .Y(n1688) );
  OAI21X1 U881 ( .A0(n5086), .A1(n1689), .B0(n1690), .Y(Inst_AEAD_u_input_n525) );
  AOI22XL U882 ( .A0(Inst_AEAD_u_input_N142), .A1(n1659), .B0(
        Inst_AEAD_u_input_sgmt_len_14_), .B1(n1660), .Y(n1690) );
  NOR3X1 U883 ( .A(n1691), .B(Inst_AEAD_u_input_n554), .C(n1660), .Y(n1659) );
  NOR2X1 U884 ( .A(Inst_AEAD_u_input_n392), .B(Inst_AEAD_u_input_n554), .Y(
        n1660) );
  OAI32XL U885 ( .A0(n1692), .A1(rst), .A2(n1693), .B0(n1694), .B1(n1657), .Y(
        Inst_AEAD_u_input_n524) );
  AOI211X1 U886 ( .A0(n1566), .A1(n1695), .B0(n1696), .C0(n1697), .Y(n1692) );
  OAI2BB1X1 U887 ( .A0N(n1698), .A1N(n1699), .B0(n1700), .Y(n1696) );
  OAI32XL U888 ( .A0(n1701), .A1(rst), .A2(n1693), .B0(n1702), .B1(n1657), .Y(
        Inst_AEAD_u_input_n523) );
  CLKNAND2X2 U889 ( .A(n1693), .B(n981), .Y(n1657) );
  CLKINVX1 U890 ( .A(n1703), .Y(n1693) );
  NOR3X1 U891 ( .A(n1697), .B(Inst_AEAD_u_input_n554), .C(n1704), .Y(n1701) );
  OAI2BB1X1 U892 ( .A0N(n1652), .A1N(Inst_AEAD_u_input_is_extra), .B0(n1705), 
        .Y(n1697) );
  AOI32XL U893 ( .A0(Inst_AEAD_u_input_n358), .A1(n468), .A2(n1706), .B0(n1695), .B1(n1619), .Y(n1705) );
  OR2X1 U894 ( .A(n1706), .B(n1652), .Y(n1695) );
  NOR2X1 U895 ( .A(rst), .B(n1707), .Y(Inst_AEAD_u_input_n522) );
  AOI31X1 U896 ( .A0(n1699), .A1(pdi_data[30]), .A2(pdi_data[28]), .B0(n1708), 
        .Y(n1707) );
  OA21X1 U897 ( .A0(n1604), .A1(n1605), .B0(Inst_AEAD_key_update), .Y(n1708)
         );
  NOR3X1 U898 ( .A(n1709), .B(pdi_data[31]), .C(n1710), .Y(n1699) );
  NOR2X1 U899 ( .A(rst), .B(n1711), .Y(Inst_AEAD_u_input_n521) );
  AOI21BX1 U900 ( .A0(Inst_AEAD_bdi_valid), .A1(n1653), .B0N(n1655), .Y(n1711)
         );
  NAND3XL U901 ( .A(n1606), .B(n1703), .C(Inst_AEAD_u_input_ctr_0_), .Y(n1655)
         );
  OAI2B11X1 U902 ( .A1N(pdi_valid), .A0(n1712), .B0(n471), .C0(n1713), .Y(
        n1703) );
  AOI21X1 U903 ( .A0(Inst_AEAD_cmd_wr_ready), .A1(Inst_AEAD_u_input_n554), 
        .B0(Inst_AEAD_u_input_n553), .Y(n1712) );
  CLKNAND2X2 U904 ( .A(Inst_AEAD_bdi_valid), .B(n1714), .Y(n1653) );
  OAI22X1 U905 ( .A0(Inst_AEAD_u_input_n321), .A1(n472), .B0(n1614), .B1(n1661), .Y(Inst_AEAD_u_input_n520) );
  OAI22X1 U906 ( .A0(Inst_AEAD_u_input_n320), .A1(n472), .B0(n1614), .B1(n1664), .Y(Inst_AEAD_u_input_n519) );
  OAI22X1 U907 ( .A0(Inst_AEAD_u_input_n319), .A1(n472), .B0(n1614), .B1(n1666), .Y(Inst_AEAD_u_input_n518) );
  OAI22X1 U908 ( .A0(Inst_AEAD_u_input_n318), .A1(n472), .B0(n1614), .B1(n1668), .Y(Inst_AEAD_u_input_n517) );
  OAI22X1 U909 ( .A0(Inst_AEAD_u_input_n317), .A1(n472), .B0(n1614), .B1(n1670), .Y(Inst_AEAD_u_input_n516) );
  OAI22X1 U910 ( .A0(Inst_AEAD_u_input_n316), .A1(n472), .B0(n1614), .B1(n1672), .Y(Inst_AEAD_u_input_n515) );
  OAI22X1 U911 ( .A0(Inst_AEAD_u_input_n315), .A1(n472), .B0(n1614), .B1(n1674), .Y(Inst_AEAD_u_input_n514) );
  OAI22X1 U912 ( .A0(Inst_AEAD_u_input_n314), .A1(n472), .B0(n1614), .B1(n1677), .Y(Inst_AEAD_u_input_n513) );
  OAI22X1 U913 ( .A0(Inst_AEAD_u_input_n313), .A1(n472), .B0(n1614), .B1(n1679), .Y(Inst_AEAD_u_input_n512) );
  OAI22X1 U914 ( .A0(Inst_AEAD_u_input_n312), .A1(n472), .B0(n1614), .B1(n1681), .Y(Inst_AEAD_u_input_n511) );
  OAI22X1 U915 ( .A0(Inst_AEAD_u_input_n311), .A1(n472), .B0(n1614), .B1(n1683), .Y(Inst_AEAD_u_input_n510) );
  OAI22X1 U916 ( .A0(Inst_AEAD_u_input_n310), .A1(n472), .B0(n1614), .B1(n1685), .Y(Inst_AEAD_u_input_n509) );
  OAI22X1 U917 ( .A0(Inst_AEAD_u_input_n309), .A1(n472), .B0(n1614), .B1(n1687), .Y(Inst_AEAD_u_input_n508) );
  OAI22X1 U918 ( .A0(Inst_AEAD_u_input_n308), .A1(n472), .B0(n1614), .B1(n1689), .Y(Inst_AEAD_u_input_n507) );
  OAI2B2X1 U919 ( .A1N(pdi_data[16]), .A0(n1614), .B0(n472), .B1(n1715), .Y(
        Inst_AEAD_u_input_n506) );
  OAI2B2X1 U920 ( .A1N(pdi_data[17]), .A0(n1614), .B0(n472), .B1(n1716), .Y(
        Inst_AEAD_u_input_n505) );
  OAI2B2X1 U921 ( .A1N(pdi_data[18]), .A0(n1614), .B0(n472), .B1(n1717), .Y(
        Inst_AEAD_u_input_n504) );
  OAI2B2X1 U922 ( .A1N(pdi_data[19]), .A0(n1614), .B0(n472), .B1(n1718), .Y(
        Inst_AEAD_u_input_n503) );
  OAI2B2X1 U923 ( .A1N(pdi_data[20]), .A0(n1614), .B0(n472), .B1(n1719), .Y(
        Inst_AEAD_u_input_n502) );
  OAI2B2X1 U924 ( .A1N(pdi_data[21]), .A0(n1614), .B0(n472), .B1(n1720), .Y(
        Inst_AEAD_u_input_n501) );
  OAI2B2X1 U925 ( .A1N(pdi_data[22]), .A0(n1614), .B0(n472), .B1(n1721), .Y(
        Inst_AEAD_u_input_n500) );
  OAI22X1 U926 ( .A0(n472), .A1(n1722), .B0(n1614), .B1(n1723), .Y(
        Inst_AEAD_u_input_n499) );
  OAI22X1 U927 ( .A0(Inst_AEAD_u_input_n307), .A1(n472), .B0(n1614), .B1(n1724), .Y(Inst_AEAD_u_input_n498) );
  OAI2B2X1 U928 ( .A1N(pdi_data[26]), .A0(n1614), .B0(n472), .B1(n1725), .Y(
        Inst_AEAD_u_input_n497) );
  OAI22X1 U929 ( .A0(n472), .A1(n1726), .B0(n1614), .B1(n1727), .Y(
        Inst_AEAD_u_input_n496) );
  OAI22X1 U930 ( .A0(Inst_AEAD_u_input_n306), .A1(n472), .B0(n1614), .B1(n1728), .Y(Inst_AEAD_u_input_n495) );
  OAI22X1 U931 ( .A0(Inst_AEAD_u_input_n305), .A1(n472), .B0(n1614), .B1(n1710), .Y(Inst_AEAD_u_input_n494) );
  OAI22X1 U932 ( .A0(Inst_AEAD_u_input_n304), .A1(n472), .B0(n1698), .B1(n1614), .Y(Inst_AEAD_u_input_n493) );
  NOR2X1 U933 ( .A(rst), .B(n1729), .Y(Inst_AEAD_u_input_n492) );
  AOI33X1 U934 ( .A0(n1730), .A1(n1709), .A2(Inst_AEAD_u_input_req_pad), .B0(
        Inst_AEAD_u_input_n554), .B1(n1731), .B2(pdi_data[25]), .Y(n1729) );
  OAI32XL U935 ( .A0(n1732), .A1(n1663), .A2(n1665), .B0(
        Inst_AEAD_u_input_n392), .B1(n1733), .Y(Inst_AEAD_u_input_n491) );
  CLKINVX1 U936 ( .A(Inst_AEAD_u_input_ploc_0_), .Y(n1733) );
  OAI32XL U937 ( .A0(n1732), .A1(Inst_AEAD_u_input_N128), .A2(n1665), .B0(
        Inst_AEAD_u_input_n392), .B1(n1734), .Y(Inst_AEAD_u_input_n490) );
  CLKINVX1 U938 ( .A(Inst_AEAD_u_input_ploc_1_), .Y(n1734) );
  OAI32XL U939 ( .A0(n1732), .A1(Inst_AEAD_u_input_sgmt_len_1_), .A2(n1663), 
        .B0(Inst_AEAD_u_input_n392), .B1(n469), .Y(Inst_AEAD_u_input_n489) );
  OAI2BB1X1 U940 ( .A0N(pdi_data[23]), .A1N(n1735), .B0(n1736), .Y(
        Inst_AEAD_u_input_n488) );
  MXI2X1 U941 ( .A(n1045), .B(Inst_AEAD_bdi[23]), .S0(n471), .Y(n1736) );
  OAI32XL U942 ( .A0(n1732), .A1(Inst_AEAD_u_input_sgmt_len_1_), .A2(
        Inst_AEAD_u_input_N128), .B0(Inst_AEAD_u_input_n392), .B1(n467), .Y(
        Inst_AEAD_u_input_n487) );
  NAND2BX1 U943 ( .AN(n1730), .B(Inst_AEAD_u_input_req_pad), .Y(n1732) );
  OAI21X1 U944 ( .A0(n1731), .A1(n1614), .B0(n1737), .Y(Inst_AEAD_u_input_n486) );
  MX2X1 U945 ( .A(Inst_AEAD_u_input_n303), .B(n467), .S0(n472), .Y(n1737) );
  CLKINVX1 U946 ( .A(n1735), .Y(n1614) );
  NOR2X1 U947 ( .A(n471), .B(Inst_AEAD_u_input_reg_sel_zero), .Y(n1735) );
  MXI2X1 U948 ( .A(Inst_AEAD_u_input_n287), .B(n1738), .S0(
        Inst_AEAD_u_input_n392), .Y(Inst_AEAD_u_input_n485) );
  AOI21X1 U949 ( .A0(Inst_AEAD_u_input_sgmt_len_1_), .A1(
        Inst_AEAD_u_input_N128), .B0(n5085), .Y(n1738) );
  MXI2X1 U950 ( .A(Inst_AEAD_u_input_n286), .B(n1739), .S0(
        Inst_AEAD_u_input_n392), .Y(Inst_AEAD_u_input_n484) );
  OAI22X1 U951 ( .A0(Inst_AEAD_u_input_n392), .A1(n1740), .B0(n1663), .B1(
        n1730), .Y(Inst_AEAD_u_input_n483) );
  OAI22X1 U952 ( .A0(Inst_AEAD_u_input_n392), .A1(n1741), .B0(n1665), .B1(
        n1730), .Y(Inst_AEAD_u_input_n482) );
  CLKNAND2X2 U953 ( .A(Inst_AEAD_u_input_n392), .B(n1691), .Y(n1730) );
  MXI2X1 U954 ( .A(n1742), .B(n1743), .S0(n1744), .Y(Inst_AEAD_u_input_n481)
         );
  CLKNAND2X2 U955 ( .A(n1745), .B(Inst_AEAD_u_input_size_0_), .Y(n1743) );
  AOI21X1 U956 ( .A0(n1745), .A1(n1740), .B0(n1746), .Y(n1742) );
  OAI22X1 U957 ( .A0(n1747), .A1(n1748), .B0(n1749), .B1(n1750), .Y(
        Inst_AEAD_u_input_n480) );
  XOR2X1 U958 ( .A(n1751), .B(n1752), .Y(n1749) );
  AOI21X1 U959 ( .A0(Inst_AEAD_u_input_size_1_), .A1(Inst_AEAD_bdi_size[1]), 
        .B0(n1753), .Y(n1752) );
  CLKNAND2X2 U960 ( .A(Inst_AEAD_u_input_size_0_), .B(Inst_AEAD_bdi_size[0]), 
        .Y(n1751) );
  OAI22X1 U961 ( .A0(n1754), .A1(n1748), .B0(n1755), .B1(n1750), .Y(
        Inst_AEAD_u_input_n479) );
  CLKINVX1 U962 ( .A(n1745), .Y(n1750) );
  XNOR2X1 U963 ( .A(n1756), .B(n1757), .Y(n1755) );
  XNOR2X1 U964 ( .A(n1567), .B(Inst_AEAD_bdi_size[2]), .Y(n1756) );
  CLKINVX1 U965 ( .A(n1746), .Y(n1748) );
  CLKINVX1 U966 ( .A(Inst_AEAD_bdi_size[2]), .Y(n1754) );
  MXI2X1 U967 ( .A(n1758), .B(n1759), .S0(Inst_AEAD_bdi_size[3]), .Y(
        Inst_AEAD_u_input_n478) );
  AOI21X1 U968 ( .A0(n1745), .A1(n1760), .B0(n1746), .Y(n1759) );
  NOR3X1 U969 ( .A(n472), .B(rst), .C(n1714), .Y(n1746) );
  NAND2BX1 U970 ( .AN(n1760), .B(n1745), .Y(n1758) );
  NOR2X1 U971 ( .A(n471), .B(rst), .Y(n1745) );
  OAI2B2X1 U972 ( .A1N(n1567), .A0(n1761), .B0(Inst_AEAD_bdi_size[2]), .B1(
        n1757), .Y(n1760) );
  AND2X1 U973 ( .A(n1757), .B(Inst_AEAD_bdi_size[2]), .Y(n1761) );
  OAI32XL U974 ( .A0(n1740), .A1(n1753), .A2(n1744), .B0(n1747), .B1(n1741), 
        .Y(n1757) );
  CLKINVX1 U975 ( .A(Inst_AEAD_u_input_size_1_), .Y(n1741) );
  CLKINVX1 U976 ( .A(Inst_AEAD_bdi_size[1]), .Y(n1747) );
  CLKINVX1 U977 ( .A(Inst_AEAD_bdi_size[0]), .Y(n1744) );
  NOR2X1 U978 ( .A(Inst_AEAD_bdi_size[1]), .B(Inst_AEAD_u_input_size_1_), .Y(
        n1753) );
  CLKINVX1 U979 ( .A(Inst_AEAD_u_input_size_0_), .Y(n1740) );
  MXI2X1 U980 ( .A(n1762), .B(n1763), .S0(n1700), .Y(Inst_AEAD_u_input_n477)
         );
  NAND3XL U981 ( .A(n1565), .B(n1764), .C(n1654), .Y(n1762) );
  AOI2BB1X1 U982 ( .A0N(n1765), .A1N(n1766), .B0(Inst_AEAD_u_input_is_extra), 
        .Y(n1654) );
  NAND3BX1 U983 ( .AN(n1767), .B(Inst_AEAD_u_input_sgmt_len_2_), .C(n1565), 
        .Y(n1766) );
  NAND4X1 U984 ( .A(n1704), .B(Inst_AEAD_u_input_n358), .C(n1663), .D(n1665), 
        .Y(n1765) );
  CLKINVX1 U985 ( .A(Inst_AEAD_u_input_sgmt_len_1_), .Y(n1665) );
  OAI31X1 U986 ( .A0(n1767), .A1(Inst_AEAD_u_input_sgmt_len_1_), .A2(
        Inst_AEAD_u_input_N128), .B0(n5085), .Y(n1764) );
  OAI2B1X1 U987 ( .A1N(Inst_AEAD_u_input_n392), .A0(n1619), .B0(n5086), .Y(
        Inst_AEAD_u_input_n421) );
  CLKINVX1 U988 ( .A(Inst_AEAD_u_input_n554), .Y(n5086) );
  CLKNAND2X2 U989 ( .A(n1739), .B(n1663), .Y(n1619) );
  CLKINVX1 U990 ( .A(Inst_AEAD_u_input_N128), .Y(n1663) );
  NOR2X1 U991 ( .A(n5085), .B(Inst_AEAD_u_input_sgmt_len_1_), .Y(n1739) );
  CLKINVX1 U992 ( .A(n1691), .Y(n5085) );
  NOR2X1 U993 ( .A(n1767), .B(Inst_AEAD_u_input_sgmt_len_2_), .Y(n1691) );
  NAND3XL U994 ( .A(n1768), .B(n1769), .C(n1770), .Y(n1767) );
  NOR4X1 U995 ( .A(n1771), .B(Inst_AEAD_u_input_sgmt_len_10_), .C(
        Inst_AEAD_u_input_sgmt_len_12_), .D(Inst_AEAD_u_input_sgmt_len_11_), 
        .Y(n1770) );
  OR3X1 U996 ( .A(Inst_AEAD_u_input_sgmt_len_14_), .B(
        Inst_AEAD_u_input_sgmt_len_15_), .C(Inst_AEAD_u_input_sgmt_len_13_), 
        .Y(n1771) );
  NOR4X1 U997 ( .A(Inst_AEAD_u_input_sgmt_len_9_), .B(
        Inst_AEAD_u_input_sgmt_len_8_), .C(Inst_AEAD_u_input_sgmt_len_7_), .D(
        Inst_AEAD_u_input_sgmt_len_6_), .Y(n1769) );
  NOR3X1 U998 ( .A(Inst_AEAD_u_input_sgmt_len_3_), .B(
        Inst_AEAD_u_input_sgmt_len_5_), .C(Inst_AEAD_u_input_sgmt_len_4_), .Y(
        n1768) );
  OAI21X1 U999 ( .A0(n1772), .A1(n1700), .B0(n1713), .Y(Inst_AEAD_u_input_n392) );
  AOI21X1 U1000 ( .A0(n1714), .A1(n1652), .B0(n1706), .Y(n1713) );
  NOR3X1 U1001 ( .A(Inst_AEAD_u_input_ps_0_), .B(Inst_AEAD_u_input_ps_2_), .C(
        n1702), .Y(n1706) );
  NOR3X1 U1002 ( .A(Inst_AEAD_u_input_ps_0_), .B(Inst_AEAD_u_input_ps_1_), .C(
        n1656), .Y(n1652) );
  CLKINVX1 U1003 ( .A(Inst_AEAD_u_input_ps_2_), .Y(n1656) );
  OAI211XL U1004 ( .A0(Inst_AEAD_u_cc_u_cc_ctrl_n52), .A1(n1773), .B0(n338), 
        .C0(n1774), .Y(n1714) );
  NOR3X1 U1005 ( .A(n868), .B(Inst_AEAD_u_cc_en_cmp), .C(n1776), .Y(n1774) );
  CLKINVX1 U1006 ( .A(n1704), .Y(n1700) );
  NOR2BX1 U1007 ( .AN(n1606), .B(Inst_AEAD_u_input_ctr_0_), .Y(n1704) );
  NOR2BX1 U1008 ( .AN(n1606), .B(n1772), .Y(Inst_AEAD_u_input_n391) );
  NOR2X1 U1009 ( .A(pdi_valid), .B(Inst_AEAD_u_input_reg_sel_zero), .Y(n1772)
         );
  NOR3X1 U1010 ( .A(n1694), .B(Inst_AEAD_u_input_ps_2_), .C(n1702), .Y(n1606)
         );
  CLKINVX1 U1011 ( .A(Inst_AEAD_u_input_ps_1_), .Y(n1702) );
  OAI221X1 U1012 ( .A0(rst), .A1(n1777), .B0(n5084), .B1(n1778), .C0(n1779), 
        .Y(Inst_AEAD_u_hdr_buffer_n435) );
  AOI22XL U1013 ( .A0(Inst_AEAD_u_hdr_buffer_n434), .A1(n1780), .B0(
        Inst_AEAD_cmd_rd_valid), .B1(Inst_AEAD_u_hdr_buffer_n431), .Y(n1779)
         );
  NOR2X1 U1014 ( .A(n1781), .B(rst), .Y(Inst_AEAD_u_hdr_buffer_n434) );
  CLKINVX1 U1015 ( .A(n1778), .Y(Inst_AEAD_u_hdr_buffer_n433) );
  CLKNAND2X2 U1016 ( .A(n1782), .B(n981), .Y(n1778) );
  OAI211XL U1017 ( .A0(Inst_AEAD_u_hdr_buffer_n374), .A1(n1781), .B0(n1783), 
        .C0(n1784), .Y(Inst_AEAD_u_hdr_buffer_n432) );
  AOI21BX1 U1018 ( .A0(n1782), .A1(n1785), .B0N(n1777), .Y(n1784) );
  AOI2BB2X1 U1019 ( .B0(n1781), .B1(Inst_AEAD_u_hdr_buffer_n374), .A0N(n1782), 
        .A1N(n1785), .Y(n1777) );
  AOI2BB1X1 U1020 ( .A0N(Inst_AEAD_u_hdr_buffer_wrptr_0_), .A1N(n1786), .B0(
        n1787), .Y(n1782) );
  AOI31X1 U1021 ( .A0(n1788), .A1(n1789), .A2(Inst_AEAD_cmd_wr_ready), .B0(rst), .Y(n1783) );
  OAI21X1 U1022 ( .A0(Inst_AEAD_u_hdr_buffer_wrptr_1_), .A1(n1787), .B0(n1788), 
        .Y(n1781) );
  OAI21BX1 U1023 ( .A0(rst), .A1(n1789), .B0N(Inst_AEAD_u_hdr_buffer_n326), 
        .Y(Inst_AEAD_u_hdr_buffer_n431) );
  MX2X1 U1024 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__23_), .B(pdi_data[31]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n430) );
  MX2X1 U1025 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__22_), .B(pdi_data[30]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n429) );
  MX2X1 U1026 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__21_), .B(pdi_data[29]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n428) );
  MX2X1 U1027 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__20_), .B(pdi_data[28]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n427) );
  MX2X1 U1028 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__19_), .B(pdi_data[27]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n426) );
  MX2X1 U1029 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__17_), .B(pdi_data[25]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n424) );
  MX2X1 U1030 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__16_), .B(pdi_data[24]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n423) );
  MX2X1 U1031 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__15_), .B(pdi_data[15]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n422) );
  MX2X1 U1032 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__14_), .B(pdi_data[14]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n421) );
  MX2X1 U1033 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__13_), .B(pdi_data[13]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n420) );
  MX2X1 U1034 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__12_), .B(pdi_data[12]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n419) );
  MX2X1 U1035 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__11_), .B(pdi_data[11]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n418) );
  MX2X1 U1036 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__10_), .B(pdi_data[10]), 
        .S0(n1612), .Y(Inst_AEAD_u_hdr_buffer_n417) );
  MX2X1 U1037 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__9_), .B(pdi_data[9]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n416) );
  MX2X1 U1038 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__8_), .B(pdi_data[8]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n415) );
  MX2X1 U1039 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__7_), .B(pdi_data[7]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n414) );
  MX2X1 U1040 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__6_), .B(pdi_data[6]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n413) );
  MX2X1 U1041 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__5_), .B(pdi_data[5]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n412) );
  MX2X1 U1042 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__4_), .B(pdi_data[4]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n411) );
  MX2X1 U1043 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__3_), .B(pdi_data[3]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n410) );
  MX2X1 U1044 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__2_), .B(pdi_data[2]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n409) );
  MX2X1 U1045 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__1_), .B(pdi_data[1]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n408) );
  MX2X1 U1046 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__0_), .B(pdi_data[0]), .S0(
        n1612), .Y(Inst_AEAD_u_hdr_buffer_n407) );
  MX2X1 U1047 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__23_), .B(pdi_data[31]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n406) );
  MX2X1 U1048 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__22_), .B(pdi_data[30]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n405) );
  MX2X1 U1049 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__21_), .B(pdi_data[29]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n404) );
  MX2X1 U1050 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__20_), .B(pdi_data[28]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n403) );
  MX2X1 U1051 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__19_), .B(pdi_data[27]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n402) );
  MX2X1 U1052 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__17_), .B(pdi_data[25]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n400) );
  MX2X1 U1053 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__16_), .B(pdi_data[24]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n399) );
  MX2X1 U1054 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__15_), .B(pdi_data[15]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n398) );
  MX2X1 U1055 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__14_), .B(pdi_data[14]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n397) );
  MX2X1 U1056 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__13_), .B(pdi_data[13]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n396) );
  MX2X1 U1057 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__12_), .B(pdi_data[12]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n395) );
  MX2X1 U1058 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__11_), .B(pdi_data[11]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n394) );
  MX2X1 U1059 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__10_), .B(pdi_data[10]), 
        .S0(n1611), .Y(Inst_AEAD_u_hdr_buffer_n393) );
  MX2X1 U1060 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__9_), .B(pdi_data[9]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n392) );
  MX2X1 U1061 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__8_), .B(pdi_data[8]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n391) );
  MX2X1 U1062 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__7_), .B(pdi_data[7]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n390) );
  MX2X1 U1063 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__6_), .B(pdi_data[6]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n389) );
  MX2X1 U1064 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__5_), .B(pdi_data[5]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n388) );
  MX2X1 U1065 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__4_), .B(pdi_data[4]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n387) );
  MX2X1 U1066 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__3_), .B(pdi_data[3]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n386) );
  MX2X1 U1067 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__2_), .B(pdi_data[2]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n385) );
  MX2X1 U1068 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__1_), .B(pdi_data[1]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n384) );
  MX2X1 U1069 ( .A(Inst_AEAD_u_hdr_buffer_memory_1__0_), .B(pdi_data[0]), .S0(
        n1611), .Y(Inst_AEAD_u_hdr_buffer_n383) );
  OAI221X1 U1070 ( .A0(n1792), .A1(n1661), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n294), .C0(n1794), .Y(
        Inst_AEAD_u_hdr_buffer_N366) );
  AOI222XL U1071 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__0_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__0_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__0_), .Y(n1794) );
  CLKINVX1 U1072 ( .A(pdi_data[0]), .Y(n1661) );
  OAI221X1 U1073 ( .A0(n1792), .A1(n1664), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n293), .C0(n1798), .Y(
        Inst_AEAD_u_hdr_buffer_N365) );
  AOI222XL U1074 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__1_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__1_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__1_), .Y(n1798) );
  CLKINVX1 U1075 ( .A(pdi_data[1]), .Y(n1664) );
  OAI221X1 U1076 ( .A0(n1792), .A1(n1666), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n292), .C0(n1799), .Y(
        Inst_AEAD_u_hdr_buffer_N364) );
  AOI222XL U1077 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__2_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__2_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__2_), .Y(n1799) );
  CLKINVX1 U1078 ( .A(pdi_data[2]), .Y(n1666) );
  OAI221X1 U1079 ( .A0(n1792), .A1(n1668), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n291), .C0(n1800), .Y(
        Inst_AEAD_u_hdr_buffer_N363) );
  AOI222XL U1080 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__3_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__3_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__3_), .Y(n1800) );
  CLKINVX1 U1081 ( .A(pdi_data[3]), .Y(n1668) );
  OAI221X1 U1082 ( .A0(n1792), .A1(n1670), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n290), .C0(n1801), .Y(
        Inst_AEAD_u_hdr_buffer_N362) );
  AOI222XL U1083 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__4_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__4_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__4_), .Y(n1801) );
  CLKINVX1 U1084 ( .A(pdi_data[4]), .Y(n1670) );
  OAI221X1 U1085 ( .A0(n1792), .A1(n1672), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n289), .C0(n1802), .Y(
        Inst_AEAD_u_hdr_buffer_N361) );
  AOI222XL U1086 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__5_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__5_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__5_), .Y(n1802) );
  CLKINVX1 U1087 ( .A(pdi_data[5]), .Y(n1672) );
  OAI221X1 U1088 ( .A0(n1792), .A1(n1674), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n288), .C0(n1803), .Y(
        Inst_AEAD_u_hdr_buffer_N360) );
  AOI222XL U1089 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__6_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__6_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__6_), .Y(n1803) );
  CLKINVX1 U1090 ( .A(pdi_data[6]), .Y(n1674) );
  OAI221X1 U1091 ( .A0(n1792), .A1(n1617), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n287), .C0(n1804), .Y(
        Inst_AEAD_u_hdr_buffer_N359) );
  AOI222XL U1092 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__7_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__7_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__7_), .Y(n1804) );
  CLKINVX1 U1093 ( .A(pdi_data[7]), .Y(n1617) );
  OAI221X1 U1094 ( .A0(n1792), .A1(n1677), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n286), .C0(n1805), .Y(
        Inst_AEAD_u_hdr_buffer_N358) );
  AOI222XL U1095 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__8_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__8_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__8_), .Y(n1805) );
  CLKINVX1 U1096 ( .A(pdi_data[8]), .Y(n1677) );
  OAI221X1 U1097 ( .A0(n1792), .A1(n1679), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n285), .C0(n1806), .Y(
        Inst_AEAD_u_hdr_buffer_N357) );
  AOI222XL U1098 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__9_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__9_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__9_), .Y(n1806) );
  CLKINVX1 U1099 ( .A(pdi_data[9]), .Y(n1679) );
  OAI221X1 U1100 ( .A0(n1792), .A1(n1681), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n284), .C0(n1807), .Y(
        Inst_AEAD_u_hdr_buffer_N356) );
  AOI222XL U1101 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__10_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__10_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__10_), .Y(n1807) );
  CLKINVX1 U1102 ( .A(pdi_data[10]), .Y(n1681) );
  OAI221X1 U1103 ( .A0(n1792), .A1(n1683), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n283), .C0(n1808), .Y(
        Inst_AEAD_u_hdr_buffer_N355) );
  AOI222XL U1104 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__11_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__11_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__11_), .Y(n1808) );
  CLKINVX1 U1105 ( .A(pdi_data[11]), .Y(n1683) );
  OAI221X1 U1106 ( .A0(n1792), .A1(n1685), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n282), .C0(n1809), .Y(
        Inst_AEAD_u_hdr_buffer_N354) );
  AOI222XL U1107 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__12_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__12_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__12_), .Y(n1809) );
  CLKINVX1 U1108 ( .A(pdi_data[12]), .Y(n1685) );
  OAI221X1 U1109 ( .A0(n1792), .A1(n1687), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n281), .C0(n1810), .Y(
        Inst_AEAD_u_hdr_buffer_N353) );
  AOI222XL U1110 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__13_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__13_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__13_), .Y(n1810) );
  CLKINVX1 U1111 ( .A(pdi_data[13]), .Y(n1687) );
  OAI221X1 U1112 ( .A0(n1792), .A1(n1689), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n280), .C0(n1811), .Y(
        Inst_AEAD_u_hdr_buffer_N352) );
  AOI222XL U1113 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__14_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__14_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__14_), .Y(n1811) );
  CLKINVX1 U1114 ( .A(pdi_data[14]), .Y(n1689) );
  OAI221X1 U1115 ( .A0(n1792), .A1(n1615), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n279), .C0(n1812), .Y(
        Inst_AEAD_u_hdr_buffer_N351) );
  AOI222XL U1116 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__15_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__15_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__15_), .Y(n1812) );
  CLKINVX1 U1117 ( .A(pdi_data[15]), .Y(n1615) );
  OAI221X1 U1118 ( .A0(n1792), .A1(n1723), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n278), .C0(n1813), .Y(
        Inst_AEAD_u_hdr_buffer_N350) );
  AOI222XL U1119 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__16_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__16_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__16_), .Y(n1813) );
  CLKINVX1 U1120 ( .A(pdi_data[24]), .Y(n1723) );
  OAI221X1 U1121 ( .A0(n1792), .A1(n1724), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n277), .C0(n1814), .Y(
        Inst_AEAD_u_hdr_buffer_N349) );
  AOI222XL U1122 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__17_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__17_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__17_), .Y(n1814) );
  CLKINVX1 U1123 ( .A(pdi_data[25]), .Y(n1724) );
  OAI221X1 U1124 ( .A0(n1613), .A1(n1815), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n276), .C0(n1816), .Y(
        Inst_AEAD_u_hdr_buffer_N348) );
  AOI22XL U1125 ( .A0(n1796), .A1(Inst_AEAD_u_hdr_buffer_memory_1__18_), .B0(
        n1797), .B1(Inst_AEAD_u_hdr_buffer_memory_0__18_), .Y(n1816) );
  CLKINVX1 U1126 ( .A(Inst_AEAD_u_hdr_buffer_memory_2__18_), .Y(n1613) );
  OAI221X1 U1127 ( .A0(n1792), .A1(n1727), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n275), .C0(n1817), .Y(
        Inst_AEAD_u_hdr_buffer_N347) );
  AOI222XL U1128 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__19_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__19_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__19_), .Y(n1817) );
  CLKINVX1 U1129 ( .A(pdi_data[27]), .Y(n1727) );
  OAI221X1 U1130 ( .A0(n1792), .A1(n1728), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n274), .C0(n1818), .Y(
        Inst_AEAD_u_hdr_buffer_N346) );
  AOI222XL U1131 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__20_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__20_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__20_), .Y(n1818) );
  CLKINVX1 U1132 ( .A(pdi_data[28]), .Y(n1728) );
  OAI221X1 U1133 ( .A0(n1792), .A1(n1710), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n273), .C0(n1819), .Y(
        Inst_AEAD_u_hdr_buffer_N345) );
  AOI222XL U1134 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__21_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__21_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__21_), .Y(n1819) );
  CLKINVX1 U1135 ( .A(pdi_data[29]), .Y(n1710) );
  OAI221X1 U1136 ( .A0(n1792), .A1(n1698), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n272), .C0(n1820), .Y(
        Inst_AEAD_u_hdr_buffer_N344) );
  AOI222XL U1137 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__22_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__22_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__22_), .Y(n1820) );
  CLKINVX1 U1138 ( .A(pdi_data[30]), .Y(n1698) );
  OAI221X1 U1139 ( .A0(n1792), .A1(n1731), .B0(n1793), .B1(
        Inst_AEAD_u_hdr_buffer_n271), .C0(n1821), .Y(
        Inst_AEAD_u_hdr_buffer_N343) );
  AOI222XL U1140 ( .A0(n1795), .A1(Inst_AEAD_u_hdr_buffer_memory_2__23_), .B0(
        n1796), .B1(Inst_AEAD_u_hdr_buffer_memory_1__23_), .C0(n1797), .C1(
        Inst_AEAD_u_hdr_buffer_memory_0__23_), .Y(n1821) );
  AND3X1 U1141 ( .A(n1610), .B(n1785), .C(n1780), .Y(n1797) );
  CLKINVX1 U1142 ( .A(n1815), .Y(n1795) );
  NAND3XL U1143 ( .A(n1785), .B(n1790), .C(Inst_AEAD_u_hdr_buffer_n374), .Y(
        n1815) );
  AOI31X1 U1144 ( .A0(n1822), .A1(n1780), .A2(n5084), .B0(n1823), .Y(n1792) );
  MX2X1 U1145 ( .A(n1824), .B(n1825), .S0(n1780), .Y(n1823) );
  NOR2X1 U1146 ( .A(n5084), .B(n1610), .Y(n1825) );
  NAND3XL U1147 ( .A(n1826), .B(n1827), .C(n1786), .Y(n1610) );
  MXI2X1 U1148 ( .A(n1788), .B(n1790), .S0(n1785), .Y(n1824) );
  NAND3XL U1149 ( .A(Inst_AEAD_u_hdr_buffer_wrptr_1_), .B(n1826), .C(n1786), 
        .Y(n1790) );
  CLKINVX1 U1150 ( .A(Inst_AEAD_u_hdr_buffer_wrptr_0_), .Y(n1826) );
  CLKINVX1 U1151 ( .A(n1791), .Y(n1822) );
  AND2X1 U1152 ( .A(n1786), .B(Inst_AEAD_u_hdr_buffer_wrptr_0_), .Y(n1787) );
  AND3X1 U1153 ( .A(pdi_valid), .B(Inst_AEAD_cmd_wr_ready), .C(n1828), .Y(
        n1786) );
  AOI32XL U1154 ( .A0(n1829), .A1(n1830), .A2(n1831), .B0(n1832), .B1(n1709), 
        .Y(n1828) );
  CLKINVX1 U1155 ( .A(Inst_AEAD_u_input_n553), .Y(n1709) );
  NOR3X1 U1156 ( .A(Inst_AEAD_u_input_ps_1_), .B(Inst_AEAD_u_input_ps_2_), .C(
        Inst_AEAD_u_input_ps_0_), .Y(Inst_AEAD_u_input_n553) );
  OAI211XL U1157 ( .A0(pdi_data[29]), .A1(n1731), .B0(Inst_AEAD_u_input_n554), 
        .C0(pdi_data[30]), .Y(n1832) );
  NOR3X1 U1158 ( .A(Inst_AEAD_u_input_ps_1_), .B(Inst_AEAD_u_input_ps_2_), .C(
        n1694), .Y(Inst_AEAD_u_input_n554) );
  CLKINVX1 U1159 ( .A(Inst_AEAD_u_input_ps_0_), .Y(n1694) );
  CLKINVX1 U1160 ( .A(pdi_data[31]), .Y(n1731) );
  XNOR2X1 U1161 ( .A(n5084), .B(Inst_AEAD_u_hdr_buffer_wrptr_0_), .Y(n1831) );
  CLKINVX1 U1162 ( .A(n1785), .Y(n5084) );
  OAI21X1 U1163 ( .A0(n1833), .A1(n376), .B0(n1834), .Y(n1785) );
  XNOR2X1 U1164 ( .A(Inst_AEAD_u_hdr_buffer_wrptr_1_), .B(
        Inst_AEAD_u_hdr_buffer_n374), .Y(n1830) );
  CLKINVX1 U1165 ( .A(n1780), .Y(Inst_AEAD_u_hdr_buffer_n374) );
  XNOR2X1 U1166 ( .A(n1834), .B(n1563), .Y(n1780) );
  CLKINVX1 U1167 ( .A(n1789), .Y(n1829) );
  OAI21X1 U1168 ( .A0(n1563), .A1(n1834), .B0(Inst_AEAD_u_hdr_buffer_looped), 
        .Y(n1789) );
  CLKNAND2X2 U1169 ( .A(n1833), .B(n376), .Y(n1834) );
  AND3X1 U1170 ( .A(Inst_AEAD_cmd_rd_ready), .B(n1835), .C(
        Inst_AEAD_cmd_rd_valid), .Y(n1833) );
  NAND3BX1 U1171 ( .AN(Inst_AEAD_u_hdr_buffer_looped), .B(n1836), .C(n1837), 
        .Y(n1835) );
  XNOR2X1 U1172 ( .A(n376), .B(Inst_AEAD_u_hdr_buffer_wrptr_0_), .Y(n1837) );
  XNOR2X1 U1173 ( .A(n1563), .B(n1827), .Y(n1836) );
  CLKINVX1 U1174 ( .A(Inst_AEAD_u_hdr_buffer_wrptr_1_), .Y(n1827) );
  CLKNAND2X2 U1175 ( .A(n1838), .B(n1621), .Y(Inst_AEAD_u_cc_u_cc_dp_n2204) );
  OR2X1 U1176 ( .A(n1839), .B(n1840), .Y(n1621) );
  MXI2X1 U1177 ( .A(n1841), .B(n1842), .S0(Inst_AEAD_u_cc_u_cc_dp_rc_2_), .Y(
        n1838) );
  AND2X1 U1178 ( .A(Inst_AEAD_u_cc_u_cc_dp_rc_1_), .B(n1622), .Y(n1841) );
  MXI2X1 U1179 ( .A(n1843), .B(n1844), .S0(Inst_AEAD_u_cc_u_cc_dp_rc_3_), .Y(
        Inst_AEAD_u_cc_u_cc_dp_n2203) );
  AOI2BB1X1 U1180 ( .A0N(n1627), .A1N(Inst_AEAD_u_cc_u_cc_dp_rc_2_), .B0(n1842), .Y(n1844) );
  OAI21BX1 U1181 ( .A0(Inst_AEAD_u_cc_u_cc_dp_rc_1_), .A1(n1627), .B0N(n1623), 
        .Y(n1842) );
  OAI21X1 U1182 ( .A0(Inst_AEAD_u_cc_u_cc_dp_rc_0_), .A1(n1627), .B0(n1625), 
        .Y(n1623) );
  NAND3XL U1183 ( .A(n1622), .B(Inst_AEAD_u_cc_u_cc_dp_rc_1_), .C(
        Inst_AEAD_u_cc_u_cc_dp_rc_2_), .Y(n1843) );
  AND3X1 U1184 ( .A(n1840), .B(n1625), .C(Inst_AEAD_u_cc_u_cc_dp_rc_0_), .Y(
        n1622) );
  CLKNAND2X2 U1185 ( .A(n1840), .B(n1845), .Y(Inst_AEAD_u_cc_u_cc_dp_n2202) );
  XNOR2X1 U1186 ( .A(n1846), .B(n1626), .Y(n1845) );
  CLKNAND2X2 U1187 ( .A(n1847), .B(n1848), .Y(Inst_AEAD_u_cc_u_cc_dp_n2201) );
  MXI2X1 U1188 ( .A(n1849), .B(n1850), .S0(Inst_AEAD_u_cc_u_cc_dp_rc_5_), .Y(
        n1847) );
  NOR3BX1 U1189 ( .AN(n1625), .B(n1627), .C(Inst_AEAD_u_cc_u_cc_dp_rc_4_), .Y(
        n1849) );
  OAI221X1 U1190 ( .A0(n1851), .A1(n377), .B0(n1627), .B1(n1852), .C0(n1848), 
        .Y(Inst_AEAD_u_cc_u_cc_dp_n2200) );
  CLKNAND2X2 U1191 ( .A(n1627), .B(n1839), .Y(n1848) );
  AOI21X1 U1192 ( .A0(Inst_AEAD_u_cc_u_cc_dp_rc_5_), .A1(n1840), .B0(n1850), 
        .Y(n1851) );
  OAI21X1 U1193 ( .A0(n1627), .A1(n1846), .B0(n1625), .Y(n1850) );
  CLKNAND2X2 U1194 ( .A(n1853), .B(n1840), .Y(Inst_AEAD_u_cc_u_cc_dp_n2199) );
  XOR2X1 U1195 ( .A(n1852), .B(Inst_AEAD_u_cc_u_cc_dp_rc_7_), .Y(n1853) );
  NAND4BX1 U1196 ( .AN(Inst_AEAD_u_cc_u_cc_dp_rc_5_), .B(n1625), .C(n1846), 
        .D(n377), .Y(n1852) );
  CLKINVX1 U1197 ( .A(Inst_AEAD_u_cc_u_cc_dp_rc_4_), .Y(n1846) );
  CLKNAND2X2 U1198 ( .A(n1626), .B(n1840), .Y(n1625) );
  OAI222X1 U1199 ( .A0(n876), .A1(n1855), .B0(n1856), .B1(n906), .C0(
        Inst_AEAD_u_input_n313), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[9]) );
  XOR2X1 U1200 ( .A(n1858), .B(n1859), .Y(n1856) );
  XOR2X1 U1201 ( .A(n1860), .B(n1861), .Y(n1858) );
  OAI222X1 U1202 ( .A0(n873), .A1(n1862), .B0(n901), .B1(n1863), .C0(n1205), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[99]) );
  XOR2X1 U1203 ( .A(n1864), .B(n1865), .Y(n1863) );
  XOR2X1 U1204 ( .A(n1866), .B(n1867), .Y(n1865) );
  OAI222X1 U1205 ( .A0(n873), .A1(n1868), .B0(n901), .B1(n1869), .C0(n1206), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[98]) );
  XOR2X1 U1206 ( .A(n1870), .B(n1871), .Y(n1869) );
  XOR2X1 U1207 ( .A(n1872), .B(n1873), .Y(n1871) );
  OAI222X1 U1208 ( .A0(n873), .A1(n1874), .B0(n901), .B1(n1875), .C0(n1207), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[97]) );
  XOR2X1 U1209 ( .A(n1876), .B(n1877), .Y(n1875) );
  XOR2X1 U1210 ( .A(n1878), .B(n1879), .Y(n1877) );
  OAI222X1 U1211 ( .A0(n873), .A1(n1880), .B0(n901), .B1(n1881), .C0(n1208), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[96]) );
  XOR2X1 U1212 ( .A(n1882), .B(n1883), .Y(n1881) );
  XOR2X1 U1213 ( .A(n1884), .B(n1885), .Y(n1883) );
  OAI222X1 U1214 ( .A0(n873), .A1(n1886), .B0(n901), .B1(n1887), .C0(n1209), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[95]) );
  XOR2X1 U1215 ( .A(n1888), .B(n1889), .Y(n1887) );
  XOR2X1 U1216 ( .A(n1890), .B(n1891), .Y(n1889) );
  OAI222X1 U1217 ( .A0(n873), .A1(n1892), .B0(n901), .B1(n1893), .C0(n1210), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[94]) );
  XOR2X1 U1218 ( .A(n1894), .B(n1895), .Y(n1893) );
  XOR2X1 U1219 ( .A(n1896), .B(n1897), .Y(n1895) );
  OAI222X1 U1220 ( .A0(n874), .A1(n1898), .B0(n901), .B1(n1899), .C0(n1211), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[93]) );
  XOR2X1 U1221 ( .A(n1900), .B(n1901), .Y(n1899) );
  XOR2X1 U1222 ( .A(n1902), .B(n1903), .Y(n1901) );
  OAI222X1 U1223 ( .A0(n873), .A1(n1904), .B0(n901), .B1(n1905), .C0(n1212), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[92]) );
  XOR2X1 U1224 ( .A(n1906), .B(n1907), .Y(n1905) );
  XOR2X1 U1225 ( .A(n1866), .B(n1908), .Y(n1907) );
  OAI222X1 U1226 ( .A0(n874), .A1(n1909), .B0(n901), .B1(n1910), .C0(n1213), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[91]) );
  XOR2X1 U1227 ( .A(n1911), .B(n1912), .Y(n1910) );
  XOR2X1 U1228 ( .A(n1872), .B(n1913), .Y(n1912) );
  OAI222X1 U1229 ( .A0(n873), .A1(n1914), .B0(n900), .B1(n1915), .C0(n1214), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[90]) );
  XOR2X1 U1230 ( .A(n1916), .B(n1917), .Y(n1915) );
  XOR2X1 U1231 ( .A(n1878), .B(n1918), .Y(n1917) );
  OAI222X1 U1232 ( .A0(n874), .A1(n1919), .B0(n1920), .B1(n906), .C0(
        Inst_AEAD_u_input_n314), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[8]) );
  XOR2X1 U1233 ( .A(n1921), .B(n1922), .Y(n1920) );
  XOR2X1 U1234 ( .A(n1923), .B(n1924), .Y(n1921) );
  OAI222X1 U1235 ( .A0(n873), .A1(n1925), .B0(n900), .B1(n1926), .C0(n1215), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[89]) );
  XOR2X1 U1236 ( .A(n1927), .B(n1928), .Y(n1926) );
  XOR2X1 U1237 ( .A(n1864), .B(n1884), .Y(n1928) );
  OAI222X1 U1238 ( .A0(n874), .A1(n1929), .B0(n900), .B1(n1930), .C0(n1216), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[88]) );
  XOR2X1 U1239 ( .A(n1931), .B(n1932), .Y(n1930) );
  XOR2X1 U1240 ( .A(n1870), .B(n1890), .Y(n1932) );
  OAI222X1 U1241 ( .A0(n873), .A1(n1933), .B0(n900), .B1(n1934), .C0(n1217), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[87]) );
  XOR2X1 U1242 ( .A(n1935), .B(n1936), .Y(n1934) );
  XOR2X1 U1243 ( .A(n1876), .B(n1896), .Y(n1936) );
  OAI222X1 U1244 ( .A0(n874), .A1(n1937), .B0(n900), .B1(n1938), .C0(n1218), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[86]) );
  XOR2X1 U1245 ( .A(n1939), .B(n1940), .Y(n1938) );
  XOR2X1 U1246 ( .A(n1882), .B(n1902), .Y(n1940) );
  OAI222X1 U1247 ( .A0(n874), .A1(n1941), .B0(n900), .B1(n1942), .C0(n1219), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[85]) );
  XOR2X1 U1248 ( .A(n1943), .B(n1944), .Y(n1942) );
  XOR2X1 U1249 ( .A(n1888), .B(n1906), .Y(n1944) );
  OAI222X1 U1250 ( .A0(n874), .A1(n1945), .B0(n900), .B1(n1946), .C0(n1220), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[84]) );
  XOR2X1 U1251 ( .A(n1947), .B(n1948), .Y(n1946) );
  XOR2X1 U1252 ( .A(n1894), .B(n1911), .Y(n1948) );
  OAI222X1 U1253 ( .A0(n874), .A1(n1949), .B0(n900), .B1(n1950), .C0(n1221), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[83]) );
  XOR2X1 U1254 ( .A(n1951), .B(n1952), .Y(n1950) );
  XOR2X1 U1255 ( .A(n1900), .B(n1916), .Y(n1952) );
  OAI222X1 U1256 ( .A0(n874), .A1(n1953), .B0(n900), .B1(n1954), .C0(n1222), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[82]) );
  XOR2X1 U1257 ( .A(n1955), .B(n1956), .Y(n1954) );
  XOR2X1 U1258 ( .A(n1864), .B(n1908), .Y(n1956) );
  XNOR2X1 U1259 ( .A(n1957), .B(n1958), .Y(n1864) );
  NOR2X1 U1260 ( .A(n1959), .B(n374), .Y(n1958) );
  OAI222X1 U1261 ( .A0(n874), .A1(n1960), .B0(n900), .B1(n1961), .C0(n1223), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[81]) );
  XOR2X1 U1262 ( .A(n1962), .B(n1963), .Y(n1961) );
  XOR2X1 U1263 ( .A(n1870), .B(n1913), .Y(n1963) );
  XNOR2X1 U1264 ( .A(n1964), .B(n1965), .Y(n1870) );
  NOR2X1 U1265 ( .A(n1966), .B(n342), .Y(n1965) );
  OAI222X1 U1266 ( .A0(n874), .A1(n1967), .B0(n900), .B1(n1968), .C0(n1224), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[80]) );
  XOR2X1 U1267 ( .A(n1969), .B(n1970), .Y(n1968) );
  XOR2X1 U1268 ( .A(n1876), .B(n1918), .Y(n1970) );
  XNOR2X1 U1269 ( .A(n1971), .B(n1972), .Y(n1876) );
  NOR2X1 U1270 ( .A(n1973), .B(n343), .Y(n1972) );
  OAI222X1 U1271 ( .A0(n874), .A1(n1974), .B0(n1975), .B1(n906), .C0(n853), 
        .C1(n1976), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[7]) );
  XOR2X1 U1272 ( .A(n1977), .B(n1978), .Y(n1975) );
  XOR2X1 U1273 ( .A(n1979), .B(n1980), .Y(n1977) );
  OAI222X1 U1274 ( .A0(n874), .A1(n1981), .B0(n899), .B1(n1982), .C0(n1225), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[79]) );
  XOR2X1 U1275 ( .A(n1983), .B(n1984), .Y(n1982) );
  XOR2X1 U1276 ( .A(n1882), .B(n1927), .Y(n1984) );
  XNOR2X1 U1277 ( .A(n1985), .B(n1986), .Y(n1882) );
  NOR2X1 U1278 ( .A(n1987), .B(n375), .Y(n1986) );
  OAI222X1 U1279 ( .A0(n874), .A1(n1988), .B0(n899), .B1(n1989), .C0(n1226), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[78]) );
  XOR2X1 U1280 ( .A(n1990), .B(n1991), .Y(n1989) );
  XOR2X1 U1281 ( .A(n1888), .B(n1931), .Y(n1991) );
  XNOR2X1 U1282 ( .A(n1992), .B(n1993), .Y(n1888) );
  AND2X1 U1283 ( .A(n1528), .B(n1994), .Y(n1993) );
  OAI222X1 U1284 ( .A0(n875), .A1(n1995), .B0(n899), .B1(n1996), .C0(n1227), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[77]) );
  XOR2X1 U1285 ( .A(n1997), .B(n1998), .Y(n1996) );
  XOR2X1 U1286 ( .A(n1894), .B(n1935), .Y(n1998) );
  XNOR2X1 U1287 ( .A(n1999), .B(n2000), .Y(n1894) );
  AND2X1 U1288 ( .A(n1527), .B(n2001), .Y(n2000) );
  OAI222X1 U1289 ( .A0(n874), .A1(n2002), .B0(n899), .B1(n2003), .C0(n1228), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[76]) );
  XOR2X1 U1290 ( .A(n2004), .B(n2005), .Y(n2003) );
  XOR2X1 U1291 ( .A(n1900), .B(n1939), .Y(n2005) );
  XNOR2X1 U1292 ( .A(n2006), .B(n2007), .Y(n1900) );
  AND2X1 U1293 ( .A(n1526), .B(n2008), .Y(n2007) );
  OAI222X1 U1294 ( .A0(n874), .A1(n2009), .B0(n899), .B1(n2010), .C0(n1229), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[75]) );
  XOR2X1 U1295 ( .A(n2011), .B(n2012), .Y(n2010) );
  XOR2X1 U1296 ( .A(n1908), .B(n1943), .Y(n2012) );
  XNOR2X1 U1297 ( .A(n2013), .B(n2014), .Y(n1908) );
  AND2X1 U1298 ( .A(n1525), .B(n2015), .Y(n2014) );
  OAI222X1 U1299 ( .A0(n874), .A1(n2016), .B0(n899), .B1(n2017), .C0(n1230), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[74]) );
  XOR2X1 U1300 ( .A(n2018), .B(n2019), .Y(n2017) );
  XOR2X1 U1301 ( .A(n1913), .B(n1947), .Y(n2019) );
  XNOR2X1 U1302 ( .A(n2020), .B(n2021), .Y(n1913) );
  AND2X1 U1303 ( .A(n1524), .B(n2022), .Y(n2021) );
  OAI222X1 U1304 ( .A0(n874), .A1(n2023), .B0(n899), .B1(n2024), .C0(n1231), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[73]) );
  XOR2X1 U1305 ( .A(n2025), .B(n2026), .Y(n2024) );
  XOR2X1 U1306 ( .A(n1918), .B(n1951), .Y(n2026) );
  XNOR2X1 U1307 ( .A(n2027), .B(n2028), .Y(n1918) );
  AND2X1 U1308 ( .A(n1523), .B(n2029), .Y(n2028) );
  OAI222X1 U1309 ( .A0(n874), .A1(n2030), .B0(n899), .B1(n2031), .C0(n1232), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[72]) );
  XOR2X1 U1310 ( .A(n2032), .B(n2033), .Y(n2031) );
  XOR2X1 U1311 ( .A(n1927), .B(n1955), .Y(n2033) );
  XNOR2X1 U1312 ( .A(n2034), .B(n2035), .Y(n1927) );
  AND2X1 U1313 ( .A(n1522), .B(n2036), .Y(n2035) );
  OAI222X1 U1314 ( .A0(n875), .A1(n2037), .B0(n899), .B1(n2038), .C0(n1233), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[71]) );
  XNOR2X1 U1315 ( .A(n2039), .B(n2040), .Y(n2038) );
  XOR2X1 U1316 ( .A(n1931), .B(n1962), .Y(n2040) );
  XNOR2X1 U1317 ( .A(n2041), .B(n2042), .Y(n1931) );
  AND2X1 U1318 ( .A(n1521), .B(n2043), .Y(n2042) );
  CLKINVX1 U1319 ( .A(n2044), .Y(n2039) );
  OAI222X1 U1320 ( .A0(n874), .A1(n2045), .B0(n899), .B1(n2046), .C0(n1234), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[70]) );
  XNOR2X1 U1321 ( .A(n2047), .B(n2048), .Y(n2046) );
  XOR2X1 U1322 ( .A(n1935), .B(n1969), .Y(n2048) );
  XNOR2X1 U1323 ( .A(n2049), .B(n2050), .Y(n1935) );
  AND2X1 U1324 ( .A(n1520), .B(n2051), .Y(n2050) );
  CLKINVX1 U1325 ( .A(n2052), .Y(n2047) );
  OAI222X1 U1326 ( .A0(n875), .A1(n2053), .B0(n2054), .B1(n907), .C0(
        Inst_AEAD_u_input_n315), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[6]) );
  XOR2X1 U1327 ( .A(n2055), .B(n2056), .Y(n2054) );
  XOR2X1 U1328 ( .A(n2057), .B(n2058), .Y(n2055) );
  OAI222X1 U1329 ( .A0(n874), .A1(n2059), .B0(n899), .B1(n2060), .C0(n1235), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[69]) );
  XNOR2X1 U1330 ( .A(n2061), .B(n2062), .Y(n2060) );
  XOR2X1 U1331 ( .A(n1939), .B(n1983), .Y(n2062) );
  XNOR2X1 U1332 ( .A(n2063), .B(n2064), .Y(n1939) );
  AND2X1 U1333 ( .A(n1519), .B(n2065), .Y(n2064) );
  CLKINVX1 U1334 ( .A(n2066), .Y(n2061) );
  OAI222X1 U1335 ( .A0(n875), .A1(n2067), .B0(n899), .B1(n2068), .C0(n1236), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[68]) );
  XNOR2X1 U1336 ( .A(n2069), .B(n2070), .Y(n2068) );
  XOR2X1 U1337 ( .A(n1943), .B(n1990), .Y(n2070) );
  XNOR2X1 U1338 ( .A(n2071), .B(n2072), .Y(n1943) );
  AND2X1 U1339 ( .A(n1518), .B(n2073), .Y(n2072) );
  CLKINVX1 U1340 ( .A(n2074), .Y(n2069) );
  OAI222X1 U1341 ( .A0(n875), .A1(n2075), .B0(n898), .B1(n2076), .C0(n1237), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[67]) );
  XNOR2X1 U1342 ( .A(n2077), .B(n2078), .Y(n2076) );
  XOR2X1 U1343 ( .A(n1947), .B(n1997), .Y(n2078) );
  XNOR2X1 U1344 ( .A(n2079), .B(n2080), .Y(n1947) );
  AND2X1 U1345 ( .A(n2081), .B(n1517), .Y(n2080) );
  CLKINVX1 U1346 ( .A(n2082), .Y(n2077) );
  OAI222X1 U1347 ( .A0(n875), .A1(n2083), .B0(n898), .B1(n2084), .C0(n1238), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[66]) );
  XNOR2X1 U1348 ( .A(n2085), .B(n2086), .Y(n2084) );
  XOR2X1 U1349 ( .A(n1951), .B(n2004), .Y(n2086) );
  XNOR2X1 U1350 ( .A(n2087), .B(n2088), .Y(n1951) );
  AND2X1 U1351 ( .A(n2089), .B(n1516), .Y(n2088) );
  CLKINVX1 U1352 ( .A(n2090), .Y(n2085) );
  OAI222X1 U1353 ( .A0(n875), .A1(n2091), .B0(n898), .B1(n2092), .C0(n1239), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[65]) );
  XNOR2X1 U1354 ( .A(n2093), .B(n2094), .Y(n2092) );
  XOR2X1 U1355 ( .A(n1955), .B(n2011), .Y(n2094) );
  XNOR2X1 U1356 ( .A(n2095), .B(n2096), .Y(n1955) );
  AND2X1 U1357 ( .A(n1515), .B(n2097), .Y(n2096) );
  CLKINVX1 U1358 ( .A(n2098), .Y(n2093) );
  OAI222X1 U1359 ( .A0(n875), .A1(n2099), .B0(n901), .B1(n2100), .C0(n1240), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[64]) );
  XNOR2X1 U1360 ( .A(n2101), .B(n2102), .Y(n2100) );
  XOR2X1 U1361 ( .A(n1962), .B(n2018), .Y(n2102) );
  XNOR2X1 U1362 ( .A(n2103), .B(n2104), .Y(n1962) );
  AND2X1 U1363 ( .A(n1514), .B(n2105), .Y(n2104) );
  OAI222X1 U1364 ( .A0(n875), .A1(n2106), .B0(n2107), .B1(n906), .C0(n1600), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[63]) );
  XOR2X1 U1365 ( .A(n2108), .B(n2109), .Y(n2107) );
  XOR2X1 U1366 ( .A(n2110), .B(n2058), .Y(n2108) );
  OAI222X1 U1367 ( .A0(n875), .A1(n2111), .B0(n2112), .B1(n905), .C0(n1568), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[62]) );
  XOR2X1 U1368 ( .A(n2113), .B(n2114), .Y(n2112) );
  XNOR2X1 U1369 ( .A(n2115), .B(n2116), .Y(n2113) );
  OAI222X1 U1370 ( .A0(n875), .A1(n2117), .B0(n2118), .B1(n907), .C0(n1569), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[61]) );
  XOR2X1 U1371 ( .A(n2119), .B(n2120), .Y(n2118) );
  XNOR2X1 U1372 ( .A(n2121), .B(n2122), .Y(n2119) );
  OAI222X1 U1373 ( .A0(n875), .A1(n2123), .B0(n2124), .B1(n905), .C0(n1570), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[60]) );
  XOR2X1 U1374 ( .A(n2125), .B(n2126), .Y(n2124) );
  XNOR2X1 U1375 ( .A(n2127), .B(n2128), .Y(n2125) );
  OAI222X1 U1376 ( .A0(n875), .A1(n2129), .B0(n2130), .B1(n906), .C0(
        Inst_AEAD_u_input_n316), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[5]) );
  XOR2X1 U1377 ( .A(n2131), .B(n2132), .Y(n2130) );
  XOR2X1 U1378 ( .A(n2133), .B(n2115), .Y(n2131) );
  OAI222X1 U1379 ( .A0(n875), .A1(n2134), .B0(n898), .B1(n2135), .C0(n1571), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[59]) );
  XOR2X1 U1380 ( .A(n2136), .B(n2137), .Y(n2135) );
  XOR2X1 U1381 ( .A(n2138), .B(n2139), .Y(n2137) );
  OAI222X1 U1382 ( .A0(n875), .A1(n2140), .B0(n898), .B1(n2141), .C0(n1572), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[58]) );
  XOR2X1 U1383 ( .A(n2142), .B(n2143), .Y(n2141) );
  XOR2X1 U1384 ( .A(n2144), .B(n2145), .Y(n2143) );
  OAI222X1 U1385 ( .A0(n875), .A1(n2146), .B0(n898), .B1(n2147), .C0(n1573), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[57]) );
  XOR2X1 U1386 ( .A(n2148), .B(n2149), .Y(n2147) );
  XOR2X1 U1387 ( .A(n2150), .B(n2151), .Y(n2149) );
  OAI222X1 U1388 ( .A0(n875), .A1(n2152), .B0(n898), .B1(n2153), .C0(n1574), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[56]) );
  XOR2X1 U1389 ( .A(n2154), .B(n2155), .Y(n2153) );
  XOR2X1 U1390 ( .A(n2156), .B(n2109), .Y(n2155) );
  OAI222X1 U1391 ( .A0(n876), .A1(n2157), .B0(n898), .B1(n2158), .C0(n1601), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[55]) );
  XOR2X1 U1392 ( .A(n2159), .B(n2160), .Y(n2158) );
  XOR2X1 U1393 ( .A(n2161), .B(n2116), .Y(n2160) );
  OAI222X1 U1394 ( .A0(n875), .A1(n2162), .B0(n898), .B1(n2163), .C0(n1575), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[54]) );
  XOR2X1 U1395 ( .A(n2164), .B(n2165), .Y(n2163) );
  XOR2X1 U1396 ( .A(n2166), .B(n2122), .Y(n2165) );
  OAI222X1 U1397 ( .A0(n876), .A1(n2167), .B0(n898), .B1(n2168), .C0(n1576), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[53]) );
  XOR2X1 U1398 ( .A(n2169), .B(n2170), .Y(n2168) );
  XOR2X1 U1399 ( .A(n2171), .B(n2128), .Y(n2170) );
  OAI222X1 U1400 ( .A0(n875), .A1(n2172), .B0(n2173), .B1(n906), .C0(n1577), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[52]) );
  XOR2X1 U1401 ( .A(n2174), .B(n2175), .Y(n2173) );
  XOR2X1 U1402 ( .A(n2176), .B(n2139), .Y(n2174) );
  OAI222X1 U1403 ( .A0(n876), .A1(n2177), .B0(n2178), .B1(n905), .C0(n1578), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[51]) );
  XOR2X1 U1404 ( .A(n2179), .B(n2180), .Y(n2178) );
  XOR2X1 U1405 ( .A(n2181), .B(n2145), .Y(n2179) );
  OAI222X1 U1406 ( .A0(n875), .A1(n2182), .B0(n897), .B1(n2183), .C0(n1579), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[50]) );
  XOR2X1 U1407 ( .A(n2184), .B(n2185), .Y(n2183) );
  XOR2X1 U1408 ( .A(n2150), .B(n1859), .Y(n2185) );
  OAI222X1 U1409 ( .A0(n876), .A1(n2186), .B0(n897), .B1(n2187), .C0(
        Inst_AEAD_u_input_n317), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[4]) );
  XOR2X1 U1410 ( .A(n2188), .B(n2189), .Y(n2187) );
  XOR2X1 U1411 ( .A(n2190), .B(n2121), .Y(n2189) );
  OAI222X1 U1412 ( .A0(n875), .A1(n2191), .B0(n897), .B1(n2192), .C0(n1580), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[49]) );
  XOR2X1 U1413 ( .A(n2193), .B(n2194), .Y(n2192) );
  XOR2X1 U1414 ( .A(n2154), .B(n1922), .Y(n2194) );
  OAI222X1 U1415 ( .A0(n876), .A1(n2195), .B0(n898), .B1(n2196), .C0(n1581), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[48]) );
  XOR2X1 U1416 ( .A(n2197), .B(n2198), .Y(n2196) );
  XOR2X1 U1417 ( .A(n2159), .B(n1978), .Y(n2198) );
  OAI222X1 U1418 ( .A0(n876), .A1(n2199), .B0(n897), .B1(n2200), .C0(n1602), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[47]) );
  XOR2X1 U1419 ( .A(n2201), .B(n2202), .Y(n2200) );
  XOR2X1 U1420 ( .A(n2164), .B(n2056), .Y(n2202) );
  OAI222X1 U1421 ( .A0(n876), .A1(n2203), .B0(n898), .B1(n2204), .C0(n1582), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[46]) );
  XOR2X1 U1422 ( .A(n2205), .B(n2206), .Y(n2204) );
  XOR2X1 U1423 ( .A(n2133), .B(n2169), .Y(n2206) );
  OAI222X1 U1424 ( .A0(n876), .A1(n2207), .B0(n2208), .B1(n906), .C0(n1583), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[45]) );
  XOR2X1 U1425 ( .A(n2209), .B(n2210), .Y(n2208) );
  XOR2X1 U1426 ( .A(n2190), .B(n2175), .Y(n2209) );
  OAI222X1 U1427 ( .A0(n876), .A1(n2211), .B0(n898), .B1(n2212), .C0(n1584), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[44]) );
  XOR2X1 U1428 ( .A(n2213), .B(n2214), .Y(n2212) );
  XOR2X1 U1429 ( .A(n2215), .B(n2180), .Y(n2214) );
  OAI222X1 U1430 ( .A0(n876), .A1(n2216), .B0(n2217), .B1(n906), .C0(n1585), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[43]) );
  XOR2X1 U1431 ( .A(n2218), .B(n2219), .Y(n2217) );
  XNOR2X1 U1432 ( .A(n2220), .B(n1859), .Y(n2218) );
  MXI2X1 U1433 ( .A(n2221), .B(n2222), .S0(n1483), .Y(n1859) );
  OAI222X1 U1434 ( .A0(n876), .A1(n2223), .B0(n2224), .B1(n905), .C0(n1586), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[42]) );
  XOR2X1 U1435 ( .A(n2225), .B(n2226), .Y(n2224) );
  XNOR2X1 U1436 ( .A(n2227), .B(n1922), .Y(n2225) );
  MXI2X1 U1437 ( .A(n2228), .B(n2229), .S0(n1482), .Y(n1922) );
  OAI222X1 U1438 ( .A0(n876), .A1(n2230), .B0(n2231), .B1(n906), .C0(n1587), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[41]) );
  XOR2X1 U1439 ( .A(n2232), .B(n2233), .Y(n2231) );
  XOR2X1 U1440 ( .A(n2234), .B(n1978), .Y(n2232) );
  MXI2X1 U1441 ( .A(n2235), .B(n2236), .S0(n1481), .Y(n1978) );
  OAI222X1 U1442 ( .A0(n876), .A1(n2237), .B0(n899), .B1(n2238), .C0(n1588), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[40]) );
  XOR2X1 U1443 ( .A(n2239), .B(n2240), .Y(n2238) );
  XOR2X1 U1444 ( .A(n2110), .B(n2056), .Y(n2240) );
  MXI2X1 U1445 ( .A(n2241), .B(n2242), .S0(n1480), .Y(n2056) );
  OAI222X1 U1446 ( .A0(n876), .A1(n2243), .B0(n2244), .B1(n906), .C0(
        Inst_AEAD_u_input_n318), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[3]) );
  XOR2X1 U1447 ( .A(n2245), .B(n2246), .Y(n2244) );
  XOR2X1 U1448 ( .A(n2215), .B(n2127), .Y(n2245) );
  OAI222X1 U1449 ( .A0(n876), .A1(n2247), .B0(n2248), .B1(n905), .C0(n1603), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[39]) );
  XOR2X1 U1450 ( .A(n2133), .B(n2249), .Y(n2248) );
  XNOR2X1 U1451 ( .A(n1860), .B(n2114), .Y(n2249) );
  MXI2X1 U1452 ( .A(n2250), .B(n2251), .S0(n1479), .Y(n2133) );
  OAI222X1 U1453 ( .A0(n876), .A1(n2252), .B0(n2253), .B1(n906), .C0(n1589), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[38]) );
  XOR2X1 U1454 ( .A(n2190), .B(n2254), .Y(n2253) );
  XNOR2X1 U1455 ( .A(n1923), .B(n2120), .Y(n2254) );
  MXI2X1 U1456 ( .A(n2255), .B(n2256), .S0(n1478), .Y(n2190) );
  OAI222X1 U1457 ( .A0(n876), .A1(n2257), .B0(n900), .B1(n2258), .C0(n1590), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[37]) );
  XOR2X1 U1458 ( .A(n2215), .B(n2259), .Y(n2258) );
  XNOR2X1 U1459 ( .A(n2126), .B(n1980), .Y(n2259) );
  MXI2X1 U1460 ( .A(n2260), .B(n2261), .S0(n1477), .Y(n2215) );
  OAI222X1 U1461 ( .A0(n876), .A1(n2262), .B0(n900), .B1(n2263), .C0(n1591), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[36]) );
  XOR2X1 U1462 ( .A(n2220), .B(n2264), .Y(n2263) );
  XOR2X1 U1463 ( .A(n2057), .B(n2136), .Y(n2264) );
  OAI222X1 U1464 ( .A0(n876), .A1(n2265), .B0(n2266), .B1(n905), .C0(n1592), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[35]) );
  XOR2X1 U1465 ( .A(n2267), .B(n2227), .Y(n2266) );
  XOR2X1 U1466 ( .A(n2142), .B(n2132), .Y(n2267) );
  OAI222X1 U1467 ( .A0(n876), .A1(n2268), .B0(n901), .B1(n2269), .C0(n1593), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[34]) );
  XOR2X1 U1468 ( .A(n2233), .B(n2270), .Y(n2269) );
  XOR2X1 U1469 ( .A(n2148), .B(n2188), .Y(n2270) );
  OAI222X1 U1470 ( .A0(n877), .A1(n2271), .B0(n897), .B1(n2272), .C0(n1594), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[33]) );
  XOR2X1 U1471 ( .A(n2246), .B(n2273), .Y(n2272) );
  XOR2X1 U1472 ( .A(n2110), .B(n2156), .Y(n2273) );
  MXI2X1 U1473 ( .A(n2274), .B(n2275), .S0(n1473), .Y(n2110) );
  OAI222X1 U1474 ( .A0(n877), .A1(n2276), .B0(n901), .B1(n2277), .C0(n1595), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[32]) );
  XOR2X1 U1475 ( .A(n2161), .B(n2278), .Y(n2277) );
  XNOR2X1 U1476 ( .A(n2114), .B(n1861), .Y(n2278) );
  MXI2X1 U1477 ( .A(n2279), .B(n2280), .S0(n1472), .Y(n2114) );
  OAI222X1 U1478 ( .A0(n877), .A1(n2281), .B0(n901), .B1(n2282), .C0(
        Inst_AEAD_u_input_n303), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[31]) );
  XOR2X1 U1479 ( .A(n2166), .B(n2283), .Y(n2282) );
  XNOR2X1 U1480 ( .A(n2120), .B(n1924), .Y(n2283) );
  MXI2X1 U1481 ( .A(n2284), .B(n2285), .S0(n1471), .Y(n2120) );
  CLKNAND2X2 U1482 ( .A(n2286), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[319]) );
  MXI2X1 U1483 ( .A(n2287), .B(n2288), .S0(n873), .Y(n2286) );
  XOR2X1 U1484 ( .A(n2289), .B(n2290), .Y(n2288) );
  XOR2X1 U1485 ( .A(n2291), .B(n2292), .Y(n2290) );
  XNOR2X1 U1486 ( .A(n1600), .B(n2293), .Y(n2287) );
  NOR2BX1 U1487 ( .AN(n2294), .B(n1560), .Y(n2293) );
  OAI222X1 U1488 ( .A0(n883), .A1(n2295), .B0(n2296), .B1(n2297), .C0(n1568), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[318]) );
  XNOR2X1 U1489 ( .A(n2298), .B(n2299), .Y(n2295) );
  XOR2X1 U1490 ( .A(n2300), .B(n2301), .Y(n2299) );
  OAI222X1 U1491 ( .A0(n883), .A1(n2302), .B0(n2303), .B1(n2297), .C0(n1569), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[317]) );
  XNOR2X1 U1492 ( .A(n2304), .B(n2305), .Y(n2302) );
  XOR2X1 U1493 ( .A(n2306), .B(n2307), .Y(n2305) );
  OAI222X1 U1494 ( .A0(n883), .A1(n2308), .B0(n2309), .B1(n2297), .C0(n1570), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[316]) );
  XNOR2X1 U1495 ( .A(n2310), .B(n2311), .Y(n2308) );
  XOR2X1 U1496 ( .A(n2312), .B(n2313), .Y(n2311) );
  OAI222X1 U1497 ( .A0(n883), .A1(n2314), .B0(n2315), .B1(n2297), .C0(n1571), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[315]) );
  XNOR2X1 U1498 ( .A(n2316), .B(n2317), .Y(n2314) );
  XOR2X1 U1499 ( .A(n2318), .B(n2319), .Y(n2317) );
  OAI222X1 U1500 ( .A0(n883), .A1(n2320), .B0(n2321), .B1(n2297), .C0(n1572), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[314]) );
  XNOR2X1 U1501 ( .A(n2322), .B(n2323), .Y(n2320) );
  XOR2X1 U1502 ( .A(n2324), .B(n2325), .Y(n2323) );
  OAI222X1 U1503 ( .A0(n883), .A1(n2326), .B0(n2327), .B1(n2297), .C0(n1573), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[313]) );
  XNOR2X1 U1504 ( .A(n2328), .B(n2329), .Y(n2326) );
  XOR2X1 U1505 ( .A(n2330), .B(n2331), .Y(n2329) );
  OAI222X1 U1506 ( .A0(n883), .A1(n2332), .B0(n2333), .B1(n2297), .C0(n1574), 
        .C1(n2294), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[312]) );
  CLKNAND2X2 U1507 ( .A(n2334), .B(n2294), .Y(n2297) );
  CLKNAND2X2 U1508 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[7]), .Y(n2294) );
  XNOR2X1 U1509 ( .A(n2336), .B(n2337), .Y(n2332) );
  XOR2X1 U1510 ( .A(n2338), .B(n2339), .Y(n2337) );
  OAI222X1 U1511 ( .A0(n883), .A1(n2340), .B0(n2341), .B1(n2342), .C0(n1601), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[311]) );
  XNOR2X1 U1512 ( .A(n2344), .B(n2345), .Y(n2340) );
  XOR2X1 U1513 ( .A(n2346), .B(n2347), .Y(n2345) );
  CLKNAND2X2 U1514 ( .A(n2348), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[310]) );
  MXI2X1 U1515 ( .A(n2349), .B(n2350), .S0(n873), .Y(n2348) );
  XOR2X1 U1516 ( .A(n2351), .B(n2352), .Y(n2350) );
  XOR2X1 U1517 ( .A(n2292), .B(n2353), .Y(n2352) );
  XNOR2X1 U1518 ( .A(n1575), .B(n2354), .Y(n2349) );
  NOR2BX1 U1519 ( .AN(n2343), .B(n1551), .Y(n2354) );
  OAI222X1 U1520 ( .A0(n877), .A1(n2355), .B0(n2356), .B1(n906), .C0(
        Inst_AEAD_u_input_n304), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[30]) );
  XOR2X1 U1521 ( .A(n2171), .B(n2357), .Y(n2356) );
  XNOR2X1 U1522 ( .A(n1979), .B(n2126), .Y(n2357) );
  MXI2X1 U1523 ( .A(n2358), .B(n2359), .S0(n1470), .Y(n2126) );
  OAI222X1 U1524 ( .A0(n883), .A1(n2360), .B0(n2361), .B1(n2342), .C0(n1576), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[309]) );
  XNOR2X1 U1525 ( .A(n2362), .B(n2363), .Y(n2360) );
  XOR2X1 U1526 ( .A(n2301), .B(n2364), .Y(n2363) );
  OAI222X1 U1527 ( .A0(n883), .A1(n2365), .B0(n2366), .B1(n2342), .C0(n1577), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[308]) );
  XNOR2X1 U1528 ( .A(n2367), .B(n2368), .Y(n2365) );
  XOR2X1 U1529 ( .A(n2307), .B(n2369), .Y(n2368) );
  OAI222X1 U1530 ( .A0(n883), .A1(n2370), .B0(n2371), .B1(n2342), .C0(n1578), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[307]) );
  XNOR2X1 U1531 ( .A(n2372), .B(n2373), .Y(n2370) );
  XOR2X1 U1532 ( .A(n2313), .B(n2374), .Y(n2373) );
  OAI222X1 U1533 ( .A0(n883), .A1(n2375), .B0(n2376), .B1(n2342), .C0(n1579), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[306]) );
  XNOR2X1 U1534 ( .A(n2377), .B(n2378), .Y(n2375) );
  XOR2X1 U1535 ( .A(n2319), .B(n2379), .Y(n2378) );
  OAI222X1 U1536 ( .A0(n884), .A1(n2380), .B0(n2381), .B1(n2342), .C0(n1580), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[305]) );
  XNOR2X1 U1537 ( .A(n2382), .B(n2383), .Y(n2380) );
  XOR2X1 U1538 ( .A(n2325), .B(n2384), .Y(n2383) );
  OAI222X1 U1539 ( .A0(n884), .A1(n2385), .B0(n2386), .B1(n2342), .C0(n1581), 
        .C1(n2343), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[304]) );
  CLKNAND2X2 U1540 ( .A(n2334), .B(n2343), .Y(n2342) );
  CLKNAND2X2 U1541 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[6]), .Y(n2343) );
  XNOR2X1 U1542 ( .A(n2387), .B(n2388), .Y(n2385) );
  XOR2X1 U1543 ( .A(n2331), .B(n2389), .Y(n2388) );
  OAI222X1 U1544 ( .A0(n884), .A1(n2390), .B0(n2391), .B1(n2392), .C0(n1602), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[303]) );
  XNOR2X1 U1545 ( .A(n2394), .B(n2395), .Y(n2390) );
  XOR2X1 U1546 ( .A(n2339), .B(n2396), .Y(n2395) );
  OAI222X1 U1547 ( .A0(n884), .A1(n2397), .B0(n2398), .B1(n2392), .C0(n1582), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[302]) );
  XNOR2X1 U1548 ( .A(n2399), .B(n2400), .Y(n2397) );
  XOR2X1 U1549 ( .A(n2347), .B(n2401), .Y(n2400) );
  OAI222X1 U1550 ( .A0(n884), .A1(n2402), .B0(n2403), .B1(n2392), .C0(n1583), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[301]) );
  XNOR2X1 U1551 ( .A(n2404), .B(n2405), .Y(n2402) );
  XOR2X1 U1552 ( .A(n2353), .B(n2406), .Y(n2405) );
  OAI222X1 U1553 ( .A0(n884), .A1(n2407), .B0(n2408), .B1(n2392), .C0(n1584), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[300]) );
  XNOR2X1 U1554 ( .A(n2409), .B(n2410), .Y(n2407) );
  XOR2X1 U1555 ( .A(n2289), .B(n2364), .Y(n2410) );
  OAI222X1 U1556 ( .A0(n877), .A1(n2411), .B0(n2412), .B1(n905), .C0(
        Inst_AEAD_u_input_n319), .C1(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[2]) );
  XOR2X1 U1557 ( .A(n2413), .B(n2220), .Y(n2412) );
  MXI2X1 U1558 ( .A(n2414), .B(n2415), .S0(n1476), .Y(n2220) );
  XOR2X1 U1559 ( .A(n2138), .B(n1861), .Y(n2413) );
  MXI2X1 U1560 ( .A(n2416), .B(n2417), .S0(n1442), .Y(n1861) );
  OAI222X1 U1561 ( .A0(n877), .A1(n2418), .B0(n902), .B1(n2419), .C0(
        Inst_AEAD_u_input_n305), .C1(n856), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[29]) );
  XOR2X1 U1562 ( .A(n2176), .B(n2420), .Y(n2419) );
  XOR2X1 U1563 ( .A(n2136), .B(n2058), .Y(n2420) );
  MXI2X1 U1564 ( .A(n2421), .B(n2422), .S0(n1439), .Y(n2058) );
  CLKINVX1 U1565 ( .A(n2423), .Y(n2422) );
  MXI2X1 U1566 ( .A(n2424), .B(n2425), .S0(n1469), .Y(n2136) );
  CLKNAND2X2 U1567 ( .A(n2426), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[299]) );
  MXI2X1 U1568 ( .A(n2427), .B(n2428), .S0(n873), .Y(n2426) );
  XNOR2X1 U1569 ( .A(n2429), .B(n2430), .Y(n2428) );
  XOR2X1 U1570 ( .A(n2298), .B(n2369), .Y(n2430) );
  XNOR2X1 U1571 ( .A(n1585), .B(n2431), .Y(n2427) );
  NOR2X1 U1572 ( .A(n2432), .B(n1540), .Y(n2431) );
  CLKNAND2X2 U1573 ( .A(n2433), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[298]) );
  MXI2X1 U1574 ( .A(n2434), .B(n2435), .S0(n873), .Y(n2433) );
  XNOR2X1 U1575 ( .A(n2436), .B(n2437), .Y(n2435) );
  XOR2X1 U1576 ( .A(n2304), .B(n2374), .Y(n2437) );
  XNOR2X1 U1577 ( .A(n1586), .B(n2438), .Y(n2434) );
  NOR2X1 U1578 ( .A(n2432), .B(n1539), .Y(n2438) );
  CLKINVX1 U1579 ( .A(n2393), .Y(n2432) );
  OAI222X1 U1580 ( .A0(n884), .A1(n2439), .B0(n2440), .B1(n2392), .C0(n1587), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[297]) );
  XNOR2X1 U1581 ( .A(n2441), .B(n2442), .Y(n2439) );
  XOR2X1 U1582 ( .A(n2310), .B(n2379), .Y(n2442) );
  OAI222X1 U1583 ( .A0(n884), .A1(n2443), .B0(n2444), .B1(n2392), .C0(n1588), 
        .C1(n2393), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[296]) );
  CLKNAND2X2 U1584 ( .A(n2334), .B(n2393), .Y(n2392) );
  CLKNAND2X2 U1585 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[5]), .Y(n2393) );
  XNOR2X1 U1586 ( .A(n2445), .B(n2446), .Y(n2443) );
  XOR2X1 U1587 ( .A(n2316), .B(n2384), .Y(n2446) );
  OAI222X1 U1588 ( .A0(n884), .A1(n2447), .B0(n2448), .B1(n2449), .C0(n1603), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[295]) );
  XNOR2X1 U1589 ( .A(n2451), .B(n2452), .Y(n2447) );
  XOR2X1 U1590 ( .A(n2322), .B(n2389), .Y(n2452) );
  OAI222X1 U1591 ( .A0(n884), .A1(n2453), .B0(n2454), .B1(n2449), .C0(n1589), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[294]) );
  XNOR2X1 U1592 ( .A(n2455), .B(n2456), .Y(n2453) );
  XOR2X1 U1593 ( .A(n2328), .B(n2396), .Y(n2456) );
  OAI222X1 U1594 ( .A0(n884), .A1(n2457), .B0(n2458), .B1(n2449), .C0(n1590), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[293]) );
  XNOR2X1 U1595 ( .A(n2459), .B(n2460), .Y(n2457) );
  XOR2X1 U1596 ( .A(n2336), .B(n2401), .Y(n2460) );
  OAI222X1 U1597 ( .A0(n884), .A1(n2461), .B0(n2462), .B1(n2449), .C0(n1591), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[292]) );
  XOR2X1 U1598 ( .A(n2463), .B(n2464), .Y(n2461) );
  XOR2X1 U1599 ( .A(n2344), .B(n2406), .Y(n2464) );
  OAI222X1 U1600 ( .A0(n885), .A1(n2465), .B0(n2466), .B1(n2449), .C0(n1592), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[291]) );
  XOR2X1 U1601 ( .A(n2467), .B(n2468), .Y(n2465) );
  XOR2X1 U1602 ( .A(n2289), .B(n2351), .Y(n2468) );
  OAI21X1 U1603 ( .A0(n2469), .A1(n2470), .B0(n2471), .Y(n2289) );
  MXI2X1 U1604 ( .A(n2472), .B(n2473), .S0(n1496), .Y(n2471) );
  NOR2BX1 U1605 ( .AN(n2469), .B(n1432), .Y(n2473) );
  CLKNAND2X2 U1606 ( .A(n2474), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[290]) );
  MXI2X1 U1607 ( .A(n2475), .B(n2476), .S0(n873), .Y(n2474) );
  XOR2X1 U1608 ( .A(n2477), .B(n2478), .Y(n2476) );
  XOR2X1 U1609 ( .A(n2298), .B(n2362), .Y(n2478) );
  OAI21X1 U1610 ( .A0(n2479), .A1(n2480), .B0(n2481), .Y(n2298) );
  MXI2X1 U1611 ( .A(n2482), .B(n2483), .S0(n1495), .Y(n2481) );
  NOR2BX1 U1612 ( .AN(n2479), .B(n1431), .Y(n2483) );
  XNOR2X1 U1613 ( .A(n1593), .B(n2484), .Y(n2475) );
  NOR2X1 U1614 ( .A(n2485), .B(n1531), .Y(n2484) );
  OAI222X1 U1615 ( .A0(n877), .A1(n2486), .B0(n902), .B1(n2487), .C0(
        Inst_AEAD_u_input_n306), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[28]) );
  XOR2X1 U1616 ( .A(n2181), .B(n2488), .Y(n2487) );
  XOR2X1 U1617 ( .A(n2142), .B(n2115), .Y(n2488) );
  MXI2X1 U1618 ( .A(n2489), .B(n2490), .S0(n1438), .Y(n2115) );
  CLKINVX1 U1619 ( .A(n2491), .Y(n2490) );
  MXI2X1 U1620 ( .A(n2492), .B(n1959), .S0(n1468), .Y(n2142) );
  CLKNAND2X2 U1621 ( .A(n2493), .B(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[289]) );
  MXI2X1 U1622 ( .A(n2494), .B(n2495), .S0(n873), .Y(n2493) );
  XOR2X1 U1623 ( .A(n2496), .B(n2497), .Y(n2495) );
  XOR2X1 U1624 ( .A(n2304), .B(n2367), .Y(n2497) );
  OAI21X1 U1625 ( .A0(n2498), .A1(n2499), .B0(n2500), .Y(n2304) );
  MXI2X1 U1626 ( .A(n2501), .B(n2502), .S0(n1494), .Y(n2500) );
  NOR2BX1 U1627 ( .AN(n2498), .B(n1430), .Y(n2502) );
  XNOR2X1 U1628 ( .A(n1594), .B(n2503), .Y(n2494) );
  NOR2X1 U1629 ( .A(n2485), .B(n1530), .Y(n2503) );
  CLKINVX1 U1630 ( .A(n2450), .Y(n2485) );
  OAI222X1 U1631 ( .A0(n885), .A1(n2504), .B0(n2505), .B1(n2449), .C0(n1595), 
        .C1(n2450), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[288]) );
  CLKNAND2X2 U1632 ( .A(n2334), .B(n2450), .Y(n2449) );
  CLKNAND2X2 U1633 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[4]), .Y(n2450) );
  XOR2X1 U1634 ( .A(n2506), .B(n2507), .Y(n2504) );
  XOR2X1 U1635 ( .A(n2310), .B(n2372), .Y(n2507) );
  OAI21X1 U1636 ( .A0(n2508), .A1(n2509), .B0(n2510), .Y(n2310) );
  MXI2X1 U1637 ( .A(n2511), .B(n2512), .S0(n1493), .Y(n2510) );
  NOR2BX1 U1638 ( .AN(n2508), .B(n1429), .Y(n2512) );
  OAI222X1 U1639 ( .A0(n885), .A1(n2513), .B0(n2514), .B1(n2515), .C0(
        Inst_AEAD_u_input_n303), .C1(n2516), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[287]) );
  XOR2X1 U1640 ( .A(n2517), .B(n2518), .Y(n2513) );
  XOR2X1 U1641 ( .A(n2316), .B(n2377), .Y(n2518) );
  OAI21X1 U1642 ( .A0(n2519), .A1(n2520), .B0(n2521), .Y(n2316) );
  MXI2X1 U1643 ( .A(n2522), .B(n2523), .S0(n1492), .Y(n2521) );
  NOR2BX1 U1644 ( .AN(n2519), .B(n1428), .Y(n2523) );
  OAI222X1 U1645 ( .A0(n885), .A1(n2524), .B0(n2514), .B1(n2525), .C0(
        Inst_AEAD_u_input_n304), .C1(n2516), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[286]) );
  XOR2X1 U1646 ( .A(n2526), .B(n2527), .Y(n2524) );
  XOR2X1 U1647 ( .A(n2322), .B(n2382), .Y(n2527) );
  OAI21X1 U1648 ( .A0(n2528), .A1(n2529), .B0(n2530), .Y(n2322) );
  MXI2X1 U1649 ( .A(n2531), .B(n2532), .S0(n1491), .Y(n2530) );
  NOR2BX1 U1650 ( .AN(n2528), .B(n1427), .Y(n2532) );
  OAI222X1 U1651 ( .A0(n885), .A1(n2533), .B0(n2514), .B1(n2534), .C0(
        Inst_AEAD_u_input_n305), .C1(n2516), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[285]) );
  XOR2X1 U1652 ( .A(n2535), .B(n2536), .Y(n2533) );
  XOR2X1 U1653 ( .A(n2328), .B(n2387), .Y(n2536) );
  OAI21X1 U1654 ( .A0(n2537), .A1(n2538), .B0(n2539), .Y(n2328) );
  MXI2X1 U1655 ( .A(n2540), .B(n2541), .S0(n1490), .Y(n2539) );
  NOR2BX1 U1656 ( .AN(n2537), .B(n1426), .Y(n2541) );
  OAI222X1 U1657 ( .A0(n885), .A1(n2542), .B0(n2514), .B1(n2543), .C0(
        Inst_AEAD_u_input_n306), .C1(n2516), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[284]) );
  XOR2X1 U1658 ( .A(n2544), .B(n2545), .Y(n2542) );
  XOR2X1 U1659 ( .A(n2336), .B(n2394), .Y(n2545) );
  OAI21X1 U1660 ( .A0(n2546), .A1(n2547), .B0(n2548), .Y(n2336) );
  MXI2X1 U1661 ( .A(n2549), .B(n2550), .S0(n1489), .Y(n2548) );
  NOR2BX1 U1662 ( .AN(n2546), .B(n1425), .Y(n2550) );
  OAI222X1 U1663 ( .A0(n885), .A1(n2551), .B0(n2514), .B1(n2552), .C0(n1726), 
        .C1(n2516), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[283]) );
  XNOR2X1 U1664 ( .A(n2399), .B(n2553), .Y(n2551) );
  XOR2X1 U1665 ( .A(n2291), .B(n2344), .Y(n2553) );
  OAI21X1 U1666 ( .A0(n2554), .A1(n2555), .B0(n2556), .Y(n2344) );
  MXI2X1 U1667 ( .A(n2557), .B(n2558), .S0(n1488), .Y(n2556) );
  NOR2BX1 U1668 ( .AN(n2554), .B(n1424), .Y(n2558) );
  OAI222X1 U1669 ( .A0(n885), .A1(n2559), .B0(n2514), .B1(n2560), .C0(n1725), 
        .C1(n2516), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[282]) );
  XNOR2X1 U1670 ( .A(n2404), .B(n2561), .Y(n2559) );
  XOR2X1 U1671 ( .A(n2300), .B(n2351), .Y(n2561) );
  OAI21X1 U1672 ( .A0(n2562), .A1(n2563), .B0(n2564), .Y(n2351) );
  MXI2X1 U1673 ( .A(n2565), .B(n2566), .S0(n1487), .Y(n2564) );
  NOR2BX1 U1674 ( .AN(n2562), .B(n1423), .Y(n2566) );
  OAI222X1 U1675 ( .A0(n885), .A1(n2567), .B0(n2514), .B1(n2568), .C0(
        Inst_AEAD_u_input_n307), .C1(n2516), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[281]) );
  XNOR2X1 U1676 ( .A(n2409), .B(n2569), .Y(n2567) );
  XOR2X1 U1677 ( .A(n2306), .B(n2362), .Y(n2569) );
  OAI21X1 U1678 ( .A0(n2570), .A1(n2571), .B0(n2572), .Y(n2362) );
  MXI2X1 U1679 ( .A(n2573), .B(n2574), .S0(n1486), .Y(n2572) );
  NOR2BX1 U1680 ( .AN(n2570), .B(n1422), .Y(n2574) );
  OAI222X1 U1681 ( .A0(n886), .A1(n2575), .B0(n2514), .B1(n2576), .C0(n1722), 
        .C1(n2516), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[280]) );
  CLKNAND2X2 U1682 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[3]), .Y(n2516) );
  OA21X1 U1683 ( .A0(n879), .A1(Inst_AEAD_bdi_valid_bytes[3]), .B0(n2577), .Y(
        n2514) );
  XNOR2X1 U1684 ( .A(n2578), .B(n2579), .Y(n2575) );
  XOR2X1 U1685 ( .A(n2312), .B(n2367), .Y(n2579) );
  OAI21X1 U1686 ( .A0(n2580), .A1(n2581), .B0(n2582), .Y(n2367) );
  MXI2X1 U1687 ( .A(n2583), .B(n2584), .S0(n1485), .Y(n2582) );
  NOR2BX1 U1688 ( .AN(n2580), .B(n1421), .Y(n2584) );
  OAI222X1 U1689 ( .A0(n877), .A1(n2585), .B0(n902), .B1(n2586), .C0(n855), 
        .C1(n1726), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[27]) );
  XOR2X1 U1690 ( .A(n2184), .B(n2587), .Y(n2586) );
  XOR2X1 U1691 ( .A(n2148), .B(n2121), .Y(n2587) );
  MXI2X1 U1692 ( .A(n2588), .B(n2589), .S0(n1437), .Y(n2121) );
  CLKINVX1 U1693 ( .A(n2590), .Y(n2589) );
  MXI2X1 U1694 ( .A(n2591), .B(n1966), .S0(n1467), .Y(n2148) );
  OAI222X1 U1695 ( .A0(n887), .A1(n2592), .B0(n2593), .B1(n2594), .C0(n2595), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[279]) );
  XNOR2X1 U1696 ( .A(n2597), .B(n2598), .Y(n2592) );
  XOR2X1 U1697 ( .A(n2318), .B(n2372), .Y(n2598) );
  OAI21X1 U1698 ( .A0(n2599), .A1(n2600), .B0(n2601), .Y(n2372) );
  MXI2X1 U1699 ( .A(n2602), .B(n2603), .S0(n1484), .Y(n2601) );
  NOR2BX1 U1700 ( .AN(n2599), .B(n1420), .Y(n2603) );
  OAI222X1 U1701 ( .A0(n887), .A1(n2604), .B0(n2593), .B1(n2605), .C0(n1721), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[278]) );
  XNOR2X1 U1702 ( .A(n2441), .B(n2606), .Y(n2604) );
  XOR2X1 U1703 ( .A(n2324), .B(n2377), .Y(n2606) );
  OAI21X1 U1704 ( .A0(n2221), .A1(n2607), .B0(n2608), .Y(n2377) );
  MXI2X1 U1705 ( .A(n2609), .B(n2610), .S0(n1483), .Y(n2608) );
  NOR2BX1 U1706 ( .AN(n2221), .B(n1419), .Y(n2610) );
  XOR2X1 U1707 ( .A(n1355), .B(n364), .Y(n2221) );
  OAI222X1 U1708 ( .A0(n887), .A1(n2611), .B0(n2593), .B1(n2612), .C0(n1720), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[277]) );
  XNOR2X1 U1709 ( .A(n2445), .B(n2613), .Y(n2611) );
  XOR2X1 U1710 ( .A(n2330), .B(n2382), .Y(n2613) );
  OAI21X1 U1711 ( .A0(n2228), .A1(n2614), .B0(n2615), .Y(n2382) );
  MXI2X1 U1712 ( .A(n2616), .B(n2617), .S0(n1482), .Y(n2615) );
  NOR2BX1 U1713 ( .AN(n2228), .B(n1418), .Y(n2617) );
  XOR2X1 U1714 ( .A(n1354), .B(n365), .Y(n2228) );
  OAI222X1 U1715 ( .A0(n887), .A1(n2618), .B0(n2593), .B1(n2619), .C0(n1719), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[276]) );
  XNOR2X1 U1716 ( .A(n2451), .B(n2620), .Y(n2618) );
  XOR2X1 U1717 ( .A(n2338), .B(n2387), .Y(n2620) );
  OAI21X1 U1718 ( .A0(n2235), .A1(n2621), .B0(n2622), .Y(n2387) );
  MXI2X1 U1719 ( .A(n2623), .B(n2624), .S0(n1481), .Y(n2622) );
  NOR2BX1 U1720 ( .AN(n2235), .B(n1417), .Y(n2624) );
  XOR2X1 U1721 ( .A(n1353), .B(n366), .Y(n2235) );
  OAI222X1 U1722 ( .A0(n887), .A1(n2625), .B0(n2593), .B1(n2626), .C0(n1718), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[275]) );
  XNOR2X1 U1723 ( .A(n2455), .B(n2627), .Y(n2625) );
  XOR2X1 U1724 ( .A(n2346), .B(n2394), .Y(n2627) );
  OAI21X1 U1725 ( .A0(n2241), .A1(n2628), .B0(n2629), .Y(n2394) );
  MXI2X1 U1726 ( .A(n2630), .B(n2631), .S0(n1480), .Y(n2629) );
  NOR2BX1 U1727 ( .AN(n2241), .B(n1416), .Y(n2631) );
  XOR2X1 U1728 ( .A(n1352), .B(n367), .Y(n2241) );
  OAI222X1 U1729 ( .A0(n887), .A1(n2632), .B0(n2593), .B1(n2633), .C0(n1717), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[274]) );
  XNOR2X1 U1730 ( .A(n2459), .B(n2634), .Y(n2632) );
  XOR2X1 U1731 ( .A(n2292), .B(n2399), .Y(n2634) );
  OAI21X1 U1732 ( .A0(n2250), .A1(n2635), .B0(n2636), .Y(n2399) );
  MXI2X1 U1733 ( .A(n2637), .B(n2638), .S0(n1479), .Y(n2636) );
  NOR2BX1 U1734 ( .AN(n2250), .B(n1415), .Y(n2638) );
  XOR2X1 U1735 ( .A(n1351), .B(n369), .Y(n2250) );
  OAI21X1 U1736 ( .A0(n2639), .A1(n2640), .B0(n2641), .Y(n2292) );
  MXI2X1 U1737 ( .A(n2097), .B(n2642), .S0(n1451), .Y(n2641) );
  NOR2BX1 U1738 ( .AN(n2639), .B(n1387), .Y(n2642) );
  OAI222X1 U1739 ( .A0(n887), .A1(n2643), .B0(n2593), .B1(n2644), .C0(n1716), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[273]) );
  XOR2X1 U1740 ( .A(n2463), .B(n2645), .Y(n2643) );
  XOR2X1 U1741 ( .A(n2301), .B(n2404), .Y(n2645) );
  OAI21X1 U1742 ( .A0(n2255), .A1(n2646), .B0(n2647), .Y(n2404) );
  MXI2X1 U1743 ( .A(n2648), .B(n2649), .S0(n1478), .Y(n2647) );
  NOR2BX1 U1744 ( .AN(n2255), .B(n1414), .Y(n2649) );
  XOR2X1 U1745 ( .A(n1350), .B(n355), .Y(n2255) );
  OAI21X1 U1746 ( .A0(n2650), .A1(n2651), .B0(n2652), .Y(n2301) );
  MXI2X1 U1747 ( .A(n2105), .B(n2653), .S0(n1450), .Y(n2652) );
  NOR2BX1 U1748 ( .AN(n2650), .B(n1386), .Y(n2653) );
  OAI222X1 U1749 ( .A0(n887), .A1(n2654), .B0(n2593), .B1(n2655), .C0(n1715), 
        .C1(n2596), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[272]) );
  CLKNAND2X2 U1750 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[2]), .Y(n2596) );
  OA21X1 U1751 ( .A0(n879), .A1(Inst_AEAD_bdi_valid_bytes[2]), .B0(n2577), .Y(
        n2593) );
  XOR2X1 U1752 ( .A(n2467), .B(n2656), .Y(n2654) );
  XOR2X1 U1753 ( .A(n2307), .B(n2409), .Y(n2656) );
  OAI21X1 U1754 ( .A0(n2260), .A1(n2657), .B0(n2658), .Y(n2409) );
  MXI2X1 U1755 ( .A(n2659), .B(n2660), .S0(n1477), .Y(n2658) );
  NOR2BX1 U1756 ( .AN(n2260), .B(n1413), .Y(n2660) );
  XOR2X1 U1757 ( .A(n1349), .B(n357), .Y(n2260) );
  OAI21X1 U1758 ( .A0(n2661), .A1(n2662), .B0(n2663), .Y(n2307) );
  MXI2X1 U1759 ( .A(n2664), .B(n2665), .S0(n1449), .Y(n2663) );
  NOR2BX1 U1760 ( .AN(n2661), .B(n1385), .Y(n2665) );
  OAI222X1 U1761 ( .A0(n887), .A1(n2666), .B0(n2667), .B1(n2668), .C0(n2669), 
        .C1(n2670), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[271]) );
  XNOR2X1 U1762 ( .A(n2477), .B(n2671), .Y(n2666) );
  XNOR2X1 U1763 ( .A(n2313), .B(n2429), .Y(n2671) );
  CLKINVX1 U1764 ( .A(n2578), .Y(n2429) );
  OAI21X1 U1765 ( .A0(n2414), .A1(n2672), .B0(n2673), .Y(n2578) );
  MXI2X1 U1766 ( .A(n2674), .B(n2675), .S0(n1476), .Y(n2673) );
  NOR2BX1 U1767 ( .AN(n2414), .B(n1412), .Y(n2675) );
  XOR2X1 U1768 ( .A(n1348), .B(n379), .Y(n2414) );
  OAI21X1 U1769 ( .A0(n2676), .A1(n2677), .B0(n2678), .Y(n2313) );
  MXI2X1 U1770 ( .A(n2679), .B(n2680), .S0(n1448), .Y(n2678) );
  NOR2BX1 U1771 ( .AN(n2676), .B(n1384), .Y(n2680) );
  OAI222X1 U1772 ( .A0(n887), .A1(n2681), .B0(n2667), .B1(n2682), .C0(
        Inst_AEAD_u_input_n308), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[270]) );
  XNOR2X1 U1773 ( .A(n2496), .B(n2683), .Y(n2681) );
  XNOR2X1 U1774 ( .A(n2319), .B(n2436), .Y(n2683) );
  CLKINVX1 U1775 ( .A(n2597), .Y(n2436) );
  OAI21X1 U1776 ( .A0(n2684), .A1(n2685), .B0(n2686), .Y(n2597) );
  MXI2X1 U1777 ( .A(n2687), .B(n2688), .S0(n1475), .Y(n2686) );
  NOR2BX1 U1778 ( .AN(n2684), .B(n1411), .Y(n2688) );
  OAI21X1 U1779 ( .A0(n2689), .A1(n2690), .B0(n2691), .Y(n2319) );
  MXI2X1 U1780 ( .A(n2692), .B(n2693), .S0(n1447), .Y(n2691) );
  NOR2BX1 U1781 ( .AN(n2689), .B(n1383), .Y(n2693) );
  OAI222X1 U1782 ( .A0(n877), .A1(n2694), .B0(n902), .B1(n2695), .C0(n853), 
        .C1(n1725), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[26]) );
  XOR2X1 U1783 ( .A(n2193), .B(n2696), .Y(n2695) );
  XOR2X1 U1784 ( .A(n2156), .B(n2127), .Y(n2696) );
  MXI2X1 U1785 ( .A(n2697), .B(n2698), .S0(n1436), .Y(n2127) );
  CLKINVX1 U1786 ( .A(n2699), .Y(n2698) );
  MXI2X1 U1787 ( .A(n2700), .B(n1973), .S0(n1466), .Y(n2156) );
  OAI222X1 U1788 ( .A0(n886), .A1(n2701), .B0(n2667), .B1(n2702), .C0(
        Inst_AEAD_u_input_n309), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[269]) );
  XOR2X1 U1789 ( .A(n2506), .B(n2703), .Y(n2701) );
  XOR2X1 U1790 ( .A(n2325), .B(n2441), .Y(n2703) );
  OAI21X1 U1791 ( .A0(n2704), .A1(n2705), .B0(n2706), .Y(n2441) );
  MXI2X1 U1792 ( .A(n2707), .B(n2708), .S0(n1474), .Y(n2706) );
  NOR2BX1 U1793 ( .AN(n2704), .B(n1410), .Y(n2708) );
  OAI21X1 U1794 ( .A0(n2709), .A1(n2710), .B0(n2711), .Y(n2325) );
  MXI2X1 U1795 ( .A(n2712), .B(n2713), .S0(n1446), .Y(n2711) );
  NOR2BX1 U1796 ( .AN(n2709), .B(n1382), .Y(n2713) );
  OAI222X1 U1797 ( .A0(n886), .A1(n2714), .B0(n2667), .B1(n2715), .C0(
        Inst_AEAD_u_input_n310), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[268]) );
  XOR2X1 U1798 ( .A(n2517), .B(n2716), .Y(n2714) );
  XOR2X1 U1799 ( .A(n2331), .B(n2445), .Y(n2716) );
  OAI21X1 U1800 ( .A0(n2274), .A1(n2717), .B0(n2718), .Y(n2445) );
  MXI2X1 U1801 ( .A(n2719), .B(n2720), .S0(n1473), .Y(n2718) );
  NOR2BX1 U1802 ( .AN(n2274), .B(n1409), .Y(n2720) );
  XOR2X1 U1803 ( .A(n1345), .B(n363), .Y(n2274) );
  OAI21X1 U1804 ( .A0(n2721), .A1(n2722), .B0(n2723), .Y(n2331) );
  MXI2X1 U1805 ( .A(n2724), .B(n2725), .S0(n1445), .Y(n2723) );
  NOR2BX1 U1806 ( .AN(n2721), .B(n1381), .Y(n2725) );
  OAI222X1 U1807 ( .A0(n886), .A1(n2726), .B0(n2667), .B1(n2727), .C0(
        Inst_AEAD_u_input_n311), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[267]) );
  XOR2X1 U1808 ( .A(n2526), .B(n2728), .Y(n2726) );
  XOR2X1 U1809 ( .A(n2339), .B(n2451), .Y(n2728) );
  OAI2BB1X1 U1810 ( .A0N(n2279), .A1N(n2729), .B0(n2730), .Y(n2451) );
  MXI2X1 U1811 ( .A(n2280), .B(n2731), .S0(n1472), .Y(n2730) );
  NOR2X1 U1812 ( .A(n1408), .B(n2279), .Y(n2731) );
  XNOR2X1 U1813 ( .A(n1344), .B(n351), .Y(n2279) );
  OAI21X1 U1814 ( .A0(n2732), .A1(n2733), .B0(n2734), .Y(n2339) );
  MXI2X1 U1815 ( .A(n2735), .B(n2736), .S0(n1444), .Y(n2734) );
  NOR2BX1 U1816 ( .AN(n2732), .B(n1380), .Y(n2736) );
  OAI222X1 U1817 ( .A0(n886), .A1(n2737), .B0(n2667), .B1(n2738), .C0(
        Inst_AEAD_u_input_n312), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[266]) );
  XOR2X1 U1818 ( .A(n2535), .B(n2739), .Y(n2737) );
  XOR2X1 U1819 ( .A(n2347), .B(n2455), .Y(n2739) );
  OAI2BB1X1 U1820 ( .A0N(n2284), .A1N(n2740), .B0(n2741), .Y(n2455) );
  MXI2X1 U1821 ( .A(n2285), .B(n2742), .S0(n1471), .Y(n2741) );
  NOR2X1 U1822 ( .A(n1407), .B(n2284), .Y(n2742) );
  XNOR2X1 U1823 ( .A(n1343), .B(n352), .Y(n2284) );
  OAI21X1 U1824 ( .A0(n2743), .A1(n2744), .B0(n2745), .Y(n2347) );
  MXI2X1 U1825 ( .A(n2746), .B(n2747), .S0(n1443), .Y(n2745) );
  NOR2BX1 U1826 ( .AN(n2743), .B(n1379), .Y(n2747) );
  OAI222X1 U1827 ( .A0(n886), .A1(n2748), .B0(n2667), .B1(n2749), .C0(
        Inst_AEAD_u_input_n313), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[265]) );
  XOR2X1 U1828 ( .A(n2544), .B(n2750), .Y(n2748) );
  XOR2X1 U1829 ( .A(n2353), .B(n2459), .Y(n2750) );
  OAI2BB1X1 U1830 ( .A0N(n2358), .A1N(n2751), .B0(n2752), .Y(n2459) );
  MXI2X1 U1831 ( .A(n2359), .B(n2753), .S0(n1470), .Y(n2752) );
  NOR2X1 U1832 ( .A(n1406), .B(n2358), .Y(n2753) );
  XNOR2X1 U1833 ( .A(n1342), .B(n353), .Y(n2358) );
  OAI21X1 U1834 ( .A0(n2416), .A1(n2754), .B0(n2755), .Y(n2353) );
  MXI2X1 U1835 ( .A(n2756), .B(n2757), .S0(n1442), .Y(n2755) );
  NOR2BX1 U1836 ( .AN(n2416), .B(n1378), .Y(n2757) );
  XOR2X1 U1837 ( .A(n1314), .B(n372), .Y(n2416) );
  OAI222X1 U1838 ( .A0(n886), .A1(n2758), .B0(n2667), .B1(n2759), .C0(
        Inst_AEAD_u_input_n314), .C1(n2670), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[264]) );
  CLKNAND2X2 U1839 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[1]), .Y(n2670) );
  OA21X1 U1840 ( .A0(n879), .A1(Inst_AEAD_bdi_valid_bytes[1]), .B0(n2577), .Y(
        n2667) );
  XOR2X1 U1841 ( .A(n2463), .B(n2760), .Y(n2758) );
  XOR2X1 U1842 ( .A(n2291), .B(n2364), .Y(n2760) );
  OAI21X1 U1843 ( .A0(n2761), .A1(n2762), .B0(n2763), .Y(n2364) );
  MXI2X1 U1844 ( .A(n2764), .B(n2765), .S0(n1441), .Y(n2763) );
  NOR2BX1 U1845 ( .AN(n2761), .B(n1377), .Y(n2765) );
  OAI21X1 U1846 ( .A0(n2766), .A1(n2767), .B0(n2768), .Y(n2291) );
  MXI2X1 U1847 ( .A(n2022), .B(n2769), .S0(n1460), .Y(n2768) );
  NOR2BX1 U1848 ( .AN(n2766), .B(n1396), .Y(n2769) );
  OA21X1 U1849 ( .A0(n2424), .A1(n2770), .B0(n2771), .Y(n2463) );
  MXI2X1 U1850 ( .A(n2772), .B(n2773), .S0(n1469), .Y(n2771) );
  NOR2BX1 U1851 ( .AN(n2424), .B(n1405), .Y(n2773) );
  XOR2X1 U1852 ( .A(n1341), .B(n368), .Y(n2424) );
  OAI222X1 U1853 ( .A0(n886), .A1(n2774), .B0(n2775), .B1(n2776), .C0(n1976), 
        .C1(n2777), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[263]) );
  XOR2X1 U1854 ( .A(n2467), .B(n2778), .Y(n2774) );
  XOR2X1 U1855 ( .A(n2300), .B(n2369), .Y(n2778) );
  OAI21X1 U1856 ( .A0(n2779), .A1(n2780), .B0(n2781), .Y(n2369) );
  MXI2X1 U1857 ( .A(n2782), .B(n2783), .S0(n341), .Y(n2781) );
  NOR2X1 U1858 ( .A(n2784), .B(n2785), .Y(n2782) );
  OAI21X1 U1859 ( .A0(n2786), .A1(n2787), .B0(n2788), .Y(n2300) );
  MXI2X1 U1860 ( .A(n2029), .B(n2789), .S0(n1459), .Y(n2788) );
  NOR2BX1 U1861 ( .AN(n2786), .B(n1395), .Y(n2789) );
  OA21X1 U1862 ( .A0(n2492), .A1(n2790), .B0(n2791), .Y(n2467) );
  MXI2X1 U1863 ( .A(n2792), .B(n2793), .S0(n1468), .Y(n2791) );
  NOR2X1 U1864 ( .A(n1404), .B(n2794), .Y(n2793) );
  CLKINVX1 U1865 ( .A(n2794), .Y(n2492) );
  XNOR2X1 U1866 ( .A(n1340), .B(n374), .Y(n2794) );
  OAI222X1 U1867 ( .A0(n886), .A1(n2795), .B0(n2775), .B1(n2796), .C0(
        Inst_AEAD_u_input_n315), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[262]) );
  XNOR2X1 U1868 ( .A(n2477), .B(n2797), .Y(n2795) );
  XOR2X1 U1869 ( .A(n2306), .B(n2374), .Y(n2797) );
  OAI21X1 U1870 ( .A0(n2421), .A1(n2798), .B0(n2799), .Y(n2374) );
  MXI2X1 U1871 ( .A(n2423), .B(n2800), .S0(n1439), .Y(n2799) );
  NOR2BX1 U1872 ( .AN(n2421), .B(n2801), .Y(n2800) );
  XNOR2X1 U1873 ( .A(n1311), .B(n1503), .Y(n2421) );
  OAI21X1 U1874 ( .A0(n2802), .A1(n2803), .B0(n2804), .Y(n2306) );
  MXI2X1 U1875 ( .A(n2036), .B(n2805), .S0(n1458), .Y(n2804) );
  NOR2BX1 U1876 ( .AN(n2802), .B(n1394), .Y(n2805) );
  OAI21X1 U1877 ( .A0(n2591), .A1(n2806), .B0(n2807), .Y(n2477) );
  MXI2X1 U1878 ( .A(n2808), .B(n2809), .S0(n1467), .Y(n2807) );
  NOR2X1 U1879 ( .A(n1403), .B(n2810), .Y(n2809) );
  CLKINVX1 U1880 ( .A(n2810), .Y(n2591) );
  XNOR2X1 U1881 ( .A(n1339), .B(n342), .Y(n2810) );
  OAI222X1 U1882 ( .A0(n886), .A1(n2811), .B0(n2775), .B1(n2812), .C0(
        Inst_AEAD_u_input_n316), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[261]) );
  XNOR2X1 U1883 ( .A(n2496), .B(n2813), .Y(n2811) );
  XOR2X1 U1884 ( .A(n2312), .B(n2379), .Y(n2813) );
  OAI21X1 U1885 ( .A0(n2489), .A1(n2814), .B0(n2815), .Y(n2379) );
  MXI2X1 U1886 ( .A(n2491), .B(n2816), .S0(n1438), .Y(n2815) );
  NOR2BX1 U1887 ( .AN(n2489), .B(n2817), .Y(n2816) );
  XNOR2X1 U1888 ( .A(n1310), .B(n1502), .Y(n2489) );
  OAI21X1 U1889 ( .A0(n2818), .A1(n2819), .B0(n2820), .Y(n2312) );
  MXI2X1 U1890 ( .A(n2043), .B(n2821), .S0(n1457), .Y(n2820) );
  NOR2BX1 U1891 ( .AN(n2818), .B(n1393), .Y(n2821) );
  OAI21X1 U1892 ( .A0(n2700), .A1(n2822), .B0(n2823), .Y(n2496) );
  MXI2X1 U1893 ( .A(n2824), .B(n2825), .S0(n1466), .Y(n2823) );
  NOR2X1 U1894 ( .A(n1402), .B(n2826), .Y(n2825) );
  CLKINVX1 U1895 ( .A(n2826), .Y(n2700) );
  XNOR2X1 U1896 ( .A(n1338), .B(n343), .Y(n2826) );
  OAI222X1 U1897 ( .A0(n886), .A1(n2827), .B0(n2775), .B1(n2828), .C0(
        Inst_AEAD_u_input_n317), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[260]) );
  XOR2X1 U1898 ( .A(n2506), .B(n2829), .Y(n2827) );
  XOR2X1 U1899 ( .A(n2318), .B(n2384), .Y(n2829) );
  OAI21X1 U1900 ( .A0(n2588), .A1(n2830), .B0(n2831), .Y(n2384) );
  MXI2X1 U1901 ( .A(n2590), .B(n2832), .S0(n1437), .Y(n2831) );
  NOR2BX1 U1902 ( .AN(n2588), .B(n2833), .Y(n2832) );
  XNOR2X1 U1903 ( .A(n1309), .B(n1501), .Y(n2588) );
  OAI21X1 U1904 ( .A0(n2834), .A1(n2835), .B0(n2836), .Y(n2318) );
  MXI2X1 U1905 ( .A(n2051), .B(n2837), .S0(n1456), .Y(n2836) );
  NOR2BX1 U1906 ( .AN(n2834), .B(n1392), .Y(n2837) );
  OA21X1 U1907 ( .A0(n2838), .A1(n2839), .B0(n2840), .Y(n2506) );
  MXI2X1 U1908 ( .A(n2841), .B(n2842), .S0(n1465), .Y(n2840) );
  NOR2X1 U1909 ( .A(n1401), .B(n2843), .Y(n2842) );
  OAI222X1 U1910 ( .A0(n877), .A1(n2844), .B0(n2845), .B1(n905), .C0(
        Inst_AEAD_u_input_n307), .C1(n853), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[25]) );
  XOR2X1 U1911 ( .A(n2197), .B(n2846), .Y(n2845) );
  XOR2X1 U1912 ( .A(n2138), .B(n2161), .Y(n2846) );
  MXI2X1 U1913 ( .A(n2838), .B(n1987), .S0(n1465), .Y(n2161) );
  CLKINVX1 U1914 ( .A(n2843), .Y(n2838) );
  XNOR2X1 U1915 ( .A(n1337), .B(n375), .Y(n2843) );
  MXI2X1 U1916 ( .A(n2847), .B(n2848), .S0(n1435), .Y(n2138) );
  CLKINVX1 U1917 ( .A(n2849), .Y(n2848) );
  OAI222X1 U1918 ( .A0(n886), .A1(n2850), .B0(n2775), .B1(n2851), .C0(
        Inst_AEAD_u_input_n318), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[259]) );
  XOR2X1 U1919 ( .A(n2517), .B(n2852), .Y(n2850) );
  XOR2X1 U1920 ( .A(n2324), .B(n2389), .Y(n2852) );
  OAI21X1 U1921 ( .A0(n2697), .A1(n2853), .B0(n2854), .Y(n2389) );
  MXI2X1 U1922 ( .A(n2699), .B(n2855), .S0(n1436), .Y(n2854) );
  NOR2BX1 U1923 ( .AN(n2697), .B(n2856), .Y(n2855) );
  XNOR2X1 U1924 ( .A(n1308), .B(n1500), .Y(n2697) );
  OAI21X1 U1925 ( .A0(n2857), .A1(n2858), .B0(n2859), .Y(n2324) );
  MXI2X1 U1926 ( .A(n2065), .B(n2860), .S0(n1455), .Y(n2859) );
  NOR2BX1 U1927 ( .AN(n2857), .B(n1391), .Y(n2860) );
  OA21X1 U1928 ( .A0(n2861), .A1(n2862), .B0(n2863), .Y(n2517) );
  MXI2X1 U1929 ( .A(n1994), .B(n2864), .S0(n1464), .Y(n2863) );
  NOR2BX1 U1930 ( .AN(n2861), .B(n1400), .Y(n2864) );
  OAI222X1 U1931 ( .A0(n885), .A1(n2865), .B0(n2775), .B1(n2866), .C0(
        Inst_AEAD_u_input_n319), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[258]) );
  XOR2X1 U1932 ( .A(n2526), .B(n2867), .Y(n2865) );
  XOR2X1 U1933 ( .A(n2330), .B(n2396), .Y(n2867) );
  OAI21X1 U1934 ( .A0(n2847), .A1(n2868), .B0(n2869), .Y(n2396) );
  MXI2X1 U1935 ( .A(n2849), .B(n2870), .S0(n1435), .Y(n2869) );
  NOR2BX1 U1936 ( .AN(n2847), .B(n2871), .Y(n2870) );
  XNOR2X1 U1937 ( .A(n1307), .B(n1499), .Y(n2847) );
  OAI21X1 U1938 ( .A0(n2872), .A1(n2873), .B0(n2874), .Y(n2330) );
  MXI2X1 U1939 ( .A(n2073), .B(n2875), .S0(n1454), .Y(n2874) );
  NOR2BX1 U1940 ( .AN(n2872), .B(n1390), .Y(n2875) );
  OA21X1 U1941 ( .A0(n2876), .A1(n2877), .B0(n2878), .Y(n2526) );
  MXI2X1 U1942 ( .A(n2001), .B(n2879), .S0(n1463), .Y(n2878) );
  NOR2BX1 U1943 ( .AN(n2876), .B(n1399), .Y(n2879) );
  OAI222X1 U1944 ( .A0(n885), .A1(n2880), .B0(n2775), .B1(n2881), .C0(
        Inst_AEAD_u_input_n320), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[257]) );
  XOR2X1 U1945 ( .A(n2535), .B(n2882), .Y(n2880) );
  XOR2X1 U1946 ( .A(n2338), .B(n2401), .Y(n2882) );
  OAI21X1 U1947 ( .A0(n2883), .A1(n2884), .B0(n2885), .Y(n2401) );
  MXI2X1 U1948 ( .A(n2886), .B(n2887), .S0(n1434), .Y(n2885) );
  NOR2BX1 U1949 ( .AN(n2883), .B(n2888), .Y(n2887) );
  OAI2BB1X1 U1950 ( .A0N(n2889), .A1N(n2890), .B0(n2891), .Y(n2338) );
  MXI2X1 U1951 ( .A(n2081), .B(n2892), .S0(n1453), .Y(n2891) );
  NOR2X1 U1952 ( .A(n1389), .B(n2889), .Y(n2892) );
  OA21X1 U1953 ( .A0(n2893), .A1(n2894), .B0(n2895), .Y(n2535) );
  MXI2X1 U1954 ( .A(n2008), .B(n2896), .S0(n1462), .Y(n2895) );
  NOR2BX1 U1955 ( .AN(n2893), .B(n1398), .Y(n2896) );
  OAI222X1 U1956 ( .A0(n885), .A1(n2897), .B0(n2775), .B1(n2898), .C0(
        Inst_AEAD_u_input_n321), .C1(n2777), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[256]) );
  CLKNAND2X2 U1957 ( .A(n2335), .B(Inst_AEAD_bdi_valid_bytes[0]), .Y(n2777) );
  OA21X1 U1958 ( .A0(n879), .A1(Inst_AEAD_bdi_valid_bytes[0]), .B0(n2577), .Y(
        n2775) );
  NAND2BX1 U1959 ( .AN(n2335), .B(n2334), .Y(n2577) );
  NOR3X1 U1960 ( .A(n2899), .B(Inst_AEAD_u_cc_u_cc_ctrl_n52), .C(n2900), .Y(
        n2335) );
  XOR2X1 U1961 ( .A(n2544), .B(n2901), .Y(n2897) );
  XOR2X1 U1962 ( .A(n2346), .B(n2406), .Y(n2901) );
  OAI21X1 U1963 ( .A0(n2902), .A1(n2903), .B0(n2904), .Y(n2406) );
  MXI2X1 U1964 ( .A(n2905), .B(n2906), .S0(n1433), .Y(n2904) );
  NOR2BX1 U1965 ( .AN(n2902), .B(n2907), .Y(n2906) );
  OAI2BB1X1 U1966 ( .A0N(n2908), .A1N(n2909), .B0(n2910), .Y(n2346) );
  MXI2X1 U1967 ( .A(n2089), .B(n2911), .S0(n1452), .Y(n2910) );
  NOR2X1 U1968 ( .A(n1388), .B(n2908), .Y(n2911) );
  OA21X1 U1969 ( .A0(n2912), .A1(n2913), .B0(n2914), .Y(n2544) );
  MXI2X1 U1970 ( .A(n2015), .B(n2915), .S0(n1461), .Y(n2914) );
  NOR2BX1 U1971 ( .AN(n2912), .B(n1397), .Y(n2915) );
  OAI222X1 U1972 ( .A0(n1496), .A1(n2916), .B0(n1052), .B1(n2917), .C0(n2918), 
        .C1(n892), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[255]) );
  XOR2X1 U1973 ( .A(n2919), .B(n2920), .Y(n2918) );
  XOR2X1 U1974 ( .A(n2921), .B(n2922), .Y(n2920) );
  AOI21X1 U1975 ( .A0(n924), .A1(n1496), .B0(n857), .Y(n2917) );
  AOI21X1 U1976 ( .A0(n1052), .A1(n927), .B0(n961), .Y(n2916) );
  OAI222X1 U1977 ( .A0(n1495), .A1(n2924), .B0(n1056), .B1(n2925), .C0(n2926), 
        .C1(n892), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[254]) );
  XOR2X1 U1978 ( .A(n2927), .B(n2928), .Y(n2926) );
  XOR2X1 U1979 ( .A(n2929), .B(n2930), .Y(n2928) );
  AOI21X1 U1980 ( .A0(n917), .A1(n1495), .B0(n857), .Y(n2925) );
  AOI21X1 U1981 ( .A0(n1056), .A1(n928), .B0(n961), .Y(n2924) );
  OAI222X1 U1982 ( .A0(n1494), .A1(n2931), .B0(n1060), .B1(n2932), .C0(n2933), 
        .C1(n892), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[253]) );
  XOR2X1 U1983 ( .A(n2934), .B(n2935), .Y(n2933) );
  XOR2X1 U1984 ( .A(n2936), .B(n2937), .Y(n2935) );
  AOI21X1 U1985 ( .A0(n917), .A1(n1494), .B0(n857), .Y(n2932) );
  AOI21X1 U1986 ( .A0(n1060), .A1(n927), .B0(n961), .Y(n2931) );
  OAI222X1 U1987 ( .A0(n1493), .A1(n2938), .B0(n1064), .B1(n2939), .C0(n2940), 
        .C1(n892), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[252]) );
  XOR2X1 U1988 ( .A(n2941), .B(n2942), .Y(n2940) );
  XOR2X1 U1989 ( .A(n2922), .B(n2943), .Y(n2942) );
  AOI21X1 U1990 ( .A0(n917), .A1(n1493), .B0(n857), .Y(n2939) );
  AOI21X1 U1991 ( .A0(n1064), .A1(n927), .B0(n961), .Y(n2938) );
  OAI222X1 U1992 ( .A0(n1492), .A1(n2944), .B0(n1068), .B1(n2945), .C0(n2946), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[251]) );
  XOR2X1 U1993 ( .A(n2947), .B(n2948), .Y(n2946) );
  XOR2X1 U1994 ( .A(n2930), .B(n2949), .Y(n2948) );
  AOI21X1 U1995 ( .A0(n917), .A1(n1492), .B0(n857), .Y(n2945) );
  AOI21X1 U1996 ( .A0(n1068), .A1(n928), .B0(n961), .Y(n2944) );
  OAI222X1 U1997 ( .A0(n1491), .A1(n2950), .B0(n1072), .B1(n2951), .C0(n2952), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[250]) );
  XOR2X1 U1998 ( .A(n2953), .B(n2954), .Y(n2952) );
  XOR2X1 U1999 ( .A(n2937), .B(n2955), .Y(n2954) );
  AOI21X1 U2000 ( .A0(n917), .A1(n1491), .B0(n857), .Y(n2951) );
  AOI21X1 U2001 ( .A0(n1072), .A1(n929), .B0(n961), .Y(n2950) );
  OAI222X1 U2002 ( .A0(n877), .A1(n2956), .B0(n2957), .B1(n906), .C0(n853), 
        .C1(n1722), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[24]) );
  XOR2X1 U2003 ( .A(n2201), .B(n2958), .Y(n2957) );
  XOR2X1 U2004 ( .A(n2144), .B(n2166), .Y(n2958) );
  MXI2X1 U2005 ( .A(n2861), .B(n2959), .S0(n1464), .Y(n2166) );
  XNOR2X1 U2006 ( .A(n1336), .B(n1528), .Y(n2861) );
  OAI222X1 U2007 ( .A0(n1490), .A1(n2960), .B0(n1076), .B1(n2961), .C0(n2962), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[249]) );
  XOR2X1 U2008 ( .A(n2963), .B(n2964), .Y(n2962) );
  XOR2X1 U2009 ( .A(n2941), .B(n2965), .Y(n2964) );
  AOI21X1 U2010 ( .A0(n917), .A1(n1490), .B0(n857), .Y(n2961) );
  AOI21X1 U2011 ( .A0(n1076), .A1(n928), .B0(n961), .Y(n2960) );
  OAI222X1 U2012 ( .A0(n1489), .A1(n2966), .B0(n1080), .B1(n2967), .C0(n2968), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[248]) );
  XOR2X1 U2013 ( .A(n2969), .B(n2970), .Y(n2968) );
  XOR2X1 U2014 ( .A(n2947), .B(n2971), .Y(n2970) );
  AOI21X1 U2015 ( .A0(n917), .A1(n1489), .B0(n858), .Y(n2967) );
  AOI21X1 U2016 ( .A0(n1080), .A1(n929), .B0(n961), .Y(n2966) );
  OAI222X1 U2017 ( .A0(n1488), .A1(n2972), .B0(n1084), .B1(n2973), .C0(n2974), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[247]) );
  XOR2X1 U2018 ( .A(n2975), .B(n2976), .Y(n2974) );
  XOR2X1 U2019 ( .A(n2953), .B(n2977), .Y(n2976) );
  AOI21X1 U2020 ( .A0(n917), .A1(n1488), .B0(n858), .Y(n2973) );
  AOI21X1 U2021 ( .A0(n1084), .A1(n928), .B0(n961), .Y(n2972) );
  OAI222X1 U2022 ( .A0(n1487), .A1(n2978), .B0(n1088), .B1(n2979), .C0(n2980), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[246]) );
  XOR2X1 U2023 ( .A(n2981), .B(n2982), .Y(n2980) );
  XOR2X1 U2024 ( .A(n2963), .B(n2983), .Y(n2982) );
  AOI21X1 U2025 ( .A0(n917), .A1(n1487), .B0(n858), .Y(n2979) );
  AOI21X1 U2026 ( .A0(n1088), .A1(n928), .B0(n961), .Y(n2978) );
  OAI222X1 U2027 ( .A0(n1486), .A1(n2984), .B0(n1092), .B1(n2985), .C0(n2986), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[245]) );
  XOR2X1 U2028 ( .A(n2987), .B(n2988), .Y(n2986) );
  XOR2X1 U2029 ( .A(n2969), .B(n2989), .Y(n2988) );
  AOI21X1 U2030 ( .A0(n917), .A1(n1486), .B0(n858), .Y(n2985) );
  AOI21X1 U2031 ( .A0(n1092), .A1(n929), .B0(n961), .Y(n2984) );
  OAI222X1 U2032 ( .A0(n1485), .A1(n2990), .B0(n1096), .B1(n2991), .C0(n2992), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[244]) );
  XOR2X1 U2033 ( .A(n2993), .B(n2994), .Y(n2992) );
  XOR2X1 U2034 ( .A(n2975), .B(n2995), .Y(n2994) );
  AOI21X1 U2035 ( .A0(n917), .A1(n1485), .B0(n858), .Y(n2991) );
  AOI21X1 U2036 ( .A0(n1096), .A1(n928), .B0(n960), .Y(n2990) );
  OAI222X1 U2037 ( .A0(n1484), .A1(n2996), .B0(n1100), .B1(n2997), .C0(n2998), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[243]) );
  XOR2X1 U2038 ( .A(n2999), .B(n3000), .Y(n2998) );
  XOR2X1 U2039 ( .A(n2981), .B(n3001), .Y(n3000) );
  AOI21X1 U2040 ( .A0(n917), .A1(n1484), .B0(n858), .Y(n2997) );
  AOI21X1 U2041 ( .A0(n1100), .A1(n930), .B0(n960), .Y(n2996) );
  OAI222X1 U2042 ( .A0(n1483), .A1(n3002), .B0(n1104), .B1(n3003), .C0(n3004), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[242]) );
  XOR2X1 U2043 ( .A(n3005), .B(n3006), .Y(n3004) );
  XOR2X1 U2044 ( .A(n2987), .B(n3007), .Y(n3006) );
  AOI21X1 U2045 ( .A0(n918), .A1(n1483), .B0(n858), .Y(n3003) );
  AOI21X1 U2046 ( .A0(n1104), .A1(n930), .B0(n960), .Y(n3002) );
  OAI222X1 U2047 ( .A0(n1482), .A1(n3008), .B0(n1108), .B1(n3009), .C0(n3010), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[241]) );
  XOR2X1 U2048 ( .A(n3011), .B(n3012), .Y(n3010) );
  XOR2X1 U2049 ( .A(n2993), .B(n3013), .Y(n3012) );
  AOI21X1 U2050 ( .A0(n918), .A1(n1482), .B0(n859), .Y(n3009) );
  AOI21X1 U2051 ( .A0(n1108), .A1(n928), .B0(n960), .Y(n3008) );
  OAI222X1 U2052 ( .A0(n1481), .A1(n3014), .B0(n1112), .B1(n3015), .C0(n3016), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[240]) );
  XOR2X1 U2053 ( .A(n3017), .B(n3018), .Y(n3016) );
  XOR2X1 U2054 ( .A(n2999), .B(n3019), .Y(n3018) );
  AOI21X1 U2055 ( .A0(n918), .A1(n1481), .B0(n859), .Y(n3015) );
  AOI21X1 U2056 ( .A0(n1112), .A1(n928), .B0(n960), .Y(n3014) );
  OAI222X1 U2057 ( .A0(n877), .A1(n3020), .B0(n3021), .B1(n905), .C0(n853), 
        .C1(n2595), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[23]) );
  XOR2X1 U2058 ( .A(n3022), .B(n2205), .Y(n3021) );
  XOR2X1 U2059 ( .A(n2171), .B(n2151), .Y(n3022) );
  MXI2X1 U2060 ( .A(n2876), .B(n3023), .S0(n1463), .Y(n2171) );
  XNOR2X1 U2061 ( .A(n1335), .B(n1527), .Y(n2876) );
  OAI222X1 U2062 ( .A0(n1480), .A1(n3024), .B0(n1116), .B1(n3025), .C0(n3026), 
        .C1(n893), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[239]) );
  XOR2X1 U2063 ( .A(n3027), .B(n3028), .Y(n3026) );
  XOR2X1 U2064 ( .A(n3005), .B(n3029), .Y(n3028) );
  AOI21X1 U2065 ( .A0(n918), .A1(n1480), .B0(n859), .Y(n3025) );
  AOI21X1 U2066 ( .A0(n1116), .A1(n929), .B0(n960), .Y(n3024) );
  OAI222X1 U2067 ( .A0(n1479), .A1(n3030), .B0(n1120), .B1(n3031), .C0(n3032), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[238]) );
  XNOR2X1 U2068 ( .A(n3033), .B(n3034), .Y(n3032) );
  XOR2X1 U2069 ( .A(n3011), .B(n3035), .Y(n3034) );
  AOI21X1 U2070 ( .A0(n918), .A1(n1479), .B0(n859), .Y(n3031) );
  AOI21X1 U2071 ( .A0(n1120), .A1(n929), .B0(n960), .Y(n3030) );
  OAI222X1 U2072 ( .A0(n1478), .A1(n3036), .B0(n1124), .B1(n3037), .C0(n3038), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[237]) );
  XNOR2X1 U2073 ( .A(n3039), .B(n3040), .Y(n3038) );
  XOR2X1 U2074 ( .A(n3017), .B(n3041), .Y(n3040) );
  AOI21X1 U2075 ( .A0(n918), .A1(n1478), .B0(n859), .Y(n3037) );
  AOI21X1 U2076 ( .A0(n1124), .A1(n929), .B0(n960), .Y(n3036) );
  OAI222X1 U2077 ( .A0(n1477), .A1(n3042), .B0(n1128), .B1(n3043), .C0(n3044), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[236]) );
  XOR2X1 U2078 ( .A(n3045), .B(n3046), .Y(n3044) );
  XOR2X1 U2079 ( .A(n3027), .B(n3047), .Y(n3046) );
  AOI21X1 U2080 ( .A0(n918), .A1(n1477), .B0(n859), .Y(n3043) );
  AOI21X1 U2081 ( .A0(n1128), .A1(n931), .B0(n960), .Y(n3042) );
  OAI222X1 U2082 ( .A0(n1476), .A1(n3048), .B0(n1132), .B1(n3049), .C0(n3050), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[235]) );
  XOR2X1 U2083 ( .A(n3051), .B(n3052), .Y(n3050) );
  XNOR2X1 U2084 ( .A(n3033), .B(n3053), .Y(n3052) );
  AOI21X1 U2085 ( .A0(n918), .A1(n1476), .B0(n859), .Y(n3049) );
  AOI21X1 U2086 ( .A0(n1132), .A1(n929), .B0(n960), .Y(n3048) );
  OAI222X1 U2087 ( .A0(n1475), .A1(n3054), .B0(n1136), .B1(n3055), .C0(n3056), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[234]) );
  XOR2X1 U2088 ( .A(n3057), .B(n3058), .Y(n3056) );
  XNOR2X1 U2089 ( .A(n3039), .B(n3059), .Y(n3058) );
  AOI21X1 U2090 ( .A0(n918), .A1(n1475), .B0(n860), .Y(n3055) );
  AOI21X1 U2091 ( .A0(n1136), .A1(n929), .B0(n960), .Y(n3054) );
  OAI222X1 U2092 ( .A0(n1474), .A1(n3060), .B0(n1140), .B1(n3061), .C0(n3062), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[233]) );
  XOR2X1 U2093 ( .A(n3063), .B(n3064), .Y(n3062) );
  XOR2X1 U2094 ( .A(n2919), .B(n3045), .Y(n3064) );
  AOI21X1 U2095 ( .A0(n918), .A1(n1474), .B0(n860), .Y(n3061) );
  AOI21X1 U2096 ( .A0(n1140), .A1(n930), .B0(n960), .Y(n3060) );
  OAI222X1 U2097 ( .A0(n1473), .A1(n3065), .B0(n1144), .B1(n3066), .C0(n3067), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[232]) );
  XOR2X1 U2098 ( .A(n3068), .B(n3069), .Y(n3067) );
  XOR2X1 U2099 ( .A(n2927), .B(n3051), .Y(n3069) );
  AOI21X1 U2100 ( .A0(n918), .A1(n1473), .B0(n860), .Y(n3066) );
  AOI21X1 U2101 ( .A0(n1144), .A1(n930), .B0(n960), .Y(n3065) );
  OAI222X1 U2102 ( .A0(n1472), .A1(n3070), .B0(n1148), .B1(n3071), .C0(n3072), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[231]) );
  XOR2X1 U2103 ( .A(n3073), .B(n3074), .Y(n3072) );
  XOR2X1 U2104 ( .A(n2934), .B(n3057), .Y(n3074) );
  AOI21X1 U2105 ( .A0(n918), .A1(n1472), .B0(n860), .Y(n3071) );
  AOI21X1 U2106 ( .A0(n1148), .A1(n930), .B0(n959), .Y(n3070) );
  OAI222X1 U2107 ( .A0(n1471), .A1(n3075), .B0(n1152), .B1(n3076), .C0(n3077), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[230]) );
  XOR2X1 U2108 ( .A(n3078), .B(n3079), .Y(n3077) );
  XOR2X1 U2109 ( .A(n2919), .B(n2943), .Y(n3079) );
  MXI2X1 U2110 ( .A(n3080), .B(n3081), .S0(n352), .Y(n2919) );
  OAI21X1 U2111 ( .A0(n1280), .A1(n3082), .B0(n3083), .Y(n3081) );
  MXI2X1 U2112 ( .A(n3084), .B(n2740), .S0(n2285), .Y(n3083) );
  OAI21X1 U2113 ( .A0(n3082), .A1(n412), .B0(n3085), .Y(n3080) );
  MXI2X1 U2114 ( .A(n2740), .B(n3084), .S0(n2285), .Y(n3085) );
  NOR2X1 U2115 ( .A(n1471), .B(n1407), .Y(n3084) );
  AND2X1 U2116 ( .A(n1407), .B(n1471), .Y(n2740) );
  AOI21X1 U2117 ( .A0(n919), .A1(n1471), .B0(n860), .Y(n3076) );
  AOI21X1 U2118 ( .A0(n1152), .A1(n930), .B0(n959), .Y(n3075) );
  OAI222X1 U2119 ( .A0(n877), .A1(n3086), .B0(n3087), .B1(n906), .C0(n853), 
        .C1(n1721), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[22]) );
  XOR2X1 U2120 ( .A(n3088), .B(n2210), .Y(n3087) );
  XOR2X1 U2121 ( .A(n2176), .B(n2109), .Y(n3088) );
  MXI2X1 U2122 ( .A(n2469), .B(n3089), .S0(n1496), .Y(n2109) );
  XNOR2X1 U2123 ( .A(n1368), .B(n1560), .Y(n2469) );
  MXI2X1 U2124 ( .A(n2893), .B(n3090), .S0(n1462), .Y(n2176) );
  XNOR2X1 U2125 ( .A(n1334), .B(n1526), .Y(n2893) );
  OAI222X1 U2126 ( .A0(n1470), .A1(n3091), .B0(n1156), .B1(n3092), .C0(n3093), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[229]) );
  XOR2X1 U2127 ( .A(n3094), .B(n3095), .Y(n3093) );
  XOR2X1 U2128 ( .A(n2927), .B(n2949), .Y(n3095) );
  MXI2X1 U2129 ( .A(n3096), .B(n3097), .S0(n353), .Y(n2927) );
  OAI21X1 U2130 ( .A0(n1279), .A1(n3098), .B0(n3099), .Y(n3097) );
  MXI2X1 U2131 ( .A(n3100), .B(n2751), .S0(n2359), .Y(n3099) );
  OAI21X1 U2132 ( .A0(n3098), .A1(n413), .B0(n3101), .Y(n3096) );
  MXI2X1 U2133 ( .A(n2751), .B(n3100), .S0(n2359), .Y(n3101) );
  NOR2X1 U2134 ( .A(n1470), .B(n1406), .Y(n3100) );
  AND2X1 U2135 ( .A(n1406), .B(n1470), .Y(n2751) );
  AOI21X1 U2136 ( .A0(n919), .A1(n1470), .B0(n860), .Y(n3092) );
  AOI21X1 U2137 ( .A0(n1156), .A1(n930), .B0(n959), .Y(n3091) );
  OAI222X1 U2138 ( .A0(n1469), .A1(n3102), .B0(n1160), .B1(n3103), .C0(n3104), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[228]) );
  XOR2X1 U2139 ( .A(n3105), .B(n3106), .Y(n3104) );
  XOR2X1 U2140 ( .A(n2934), .B(n2955), .Y(n3106) );
  MXI2X1 U2141 ( .A(n3107), .B(n3108), .S0(n368), .Y(n2934) );
  OAI21X1 U2142 ( .A0(n1278), .A1(n3109), .B0(n3110), .Y(n3108) );
  MXI2X1 U2143 ( .A(n3111), .B(n3112), .S0(n2772), .Y(n3110) );
  OAI21X1 U2144 ( .A0(n3109), .A1(n405), .B0(n3113), .Y(n3107) );
  MXI2X1 U2145 ( .A(n3112), .B(n3111), .S0(n2772), .Y(n3113) );
  CLKINVX1 U2146 ( .A(n2425), .Y(n2772) );
  NOR2X1 U2147 ( .A(n1469), .B(n1405), .Y(n3111) );
  CLKINVX1 U2148 ( .A(n2770), .Y(n3112) );
  CLKNAND2X2 U2149 ( .A(n1405), .B(n1469), .Y(n2770) );
  AOI21X1 U2150 ( .A0(n919), .A1(n1469), .B0(n860), .Y(n3103) );
  AOI21X1 U2151 ( .A0(n1160), .A1(n930), .B0(n959), .Y(n3102) );
  OAI222X1 U2152 ( .A0(n1468), .A1(n3114), .B0(n1164), .B1(n3115), .C0(n3116), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[227]) );
  XOR2X1 U2153 ( .A(n3117), .B(n3118), .Y(n3116) );
  XOR2X1 U2154 ( .A(n2943), .B(n2965), .Y(n3118) );
  MXI2X1 U2155 ( .A(n3119), .B(n3120), .S0(n374), .Y(n2943) );
  OAI21X1 U2156 ( .A0(n1277), .A1(n1957), .B0(n3121), .Y(n3120) );
  MXI2X1 U2157 ( .A(n3122), .B(n3123), .S0(n2792), .Y(n3121) );
  OAI21X1 U2158 ( .A0(n1957), .A1(n414), .B0(n3124), .Y(n3119) );
  MXI2X1 U2159 ( .A(n3123), .B(n3122), .S0(n2792), .Y(n3124) );
  CLKINVX1 U2160 ( .A(n1959), .Y(n2792) );
  XNOR2X1 U2161 ( .A(n1277), .B(n445), .Y(n1959) );
  NOR2X1 U2162 ( .A(n1468), .B(n1404), .Y(n3122) );
  CLKINVX1 U2163 ( .A(n2790), .Y(n3123) );
  CLKNAND2X2 U2164 ( .A(n1404), .B(n1468), .Y(n2790) );
  CLKINVX1 U2165 ( .A(n3125), .Y(n1957) );
  AOI21X1 U2166 ( .A0(n919), .A1(n1468), .B0(n861), .Y(n3115) );
  AOI21X1 U2167 ( .A0(n1164), .A1(n931), .B0(n959), .Y(n3114) );
  OAI222X1 U2168 ( .A0(n1467), .A1(n3126), .B0(n1168), .B1(n3127), .C0(n3128), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[226]) );
  XOR2X1 U2169 ( .A(n3129), .B(n3130), .Y(n3128) );
  XOR2X1 U2170 ( .A(n2949), .B(n2971), .Y(n3130) );
  MXI2X1 U2171 ( .A(n3131), .B(n3132), .S0(n342), .Y(n2949) );
  OAI21X1 U2172 ( .A0(n1276), .A1(n1964), .B0(n3133), .Y(n3132) );
  MXI2X1 U2173 ( .A(n3134), .B(n3135), .S0(n2808), .Y(n3133) );
  OAI21X1 U2174 ( .A0(n1964), .A1(n415), .B0(n3136), .Y(n3131) );
  MXI2X1 U2175 ( .A(n3135), .B(n3134), .S0(n2808), .Y(n3136) );
  CLKINVX1 U2176 ( .A(n1966), .Y(n2808) );
  XNOR2X1 U2177 ( .A(n1276), .B(n446), .Y(n1966) );
  NOR2X1 U2178 ( .A(n1467), .B(n1403), .Y(n3134) );
  CLKINVX1 U2179 ( .A(n2806), .Y(n3135) );
  CLKNAND2X2 U2180 ( .A(n1403), .B(n1467), .Y(n2806) );
  CLKINVX1 U2181 ( .A(n3137), .Y(n1964) );
  AOI21X1 U2182 ( .A0(n919), .A1(n1467), .B0(n861), .Y(n3127) );
  AOI21X1 U2183 ( .A0(n1168), .A1(n930), .B0(n959), .Y(n3126) );
  OAI222X1 U2184 ( .A0(n1466), .A1(n3138), .B0(n1172), .B1(n3139), .C0(n3140), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[225]) );
  XOR2X1 U2185 ( .A(n3141), .B(n3142), .Y(n3140) );
  XOR2X1 U2186 ( .A(n2955), .B(n2977), .Y(n3142) );
  MXI2X1 U2187 ( .A(n3143), .B(n3144), .S0(n343), .Y(n2955) );
  OAI21X1 U2188 ( .A0(n1275), .A1(n1971), .B0(n3145), .Y(n3144) );
  MXI2X1 U2189 ( .A(n3146), .B(n3147), .S0(n2824), .Y(n3145) );
  OAI21X1 U2190 ( .A0(n1971), .A1(n416), .B0(n3148), .Y(n3143) );
  MXI2X1 U2191 ( .A(n3147), .B(n3146), .S0(n2824), .Y(n3148) );
  CLKINVX1 U2192 ( .A(n1973), .Y(n2824) );
  XNOR2X1 U2193 ( .A(n1275), .B(n447), .Y(n1973) );
  NOR2X1 U2194 ( .A(n1466), .B(n1402), .Y(n3146) );
  CLKINVX1 U2195 ( .A(n2822), .Y(n3147) );
  CLKNAND2X2 U2196 ( .A(n1402), .B(n1466), .Y(n2822) );
  CLKINVX1 U2197 ( .A(n3149), .Y(n1971) );
  AOI21X1 U2198 ( .A0(n919), .A1(n1466), .B0(n861), .Y(n3139) );
  AOI21X1 U2199 ( .A0(n1172), .A1(n931), .B0(n959), .Y(n3138) );
  OAI222X1 U2200 ( .A0(n1465), .A1(n3150), .B0(n1176), .B1(n3151), .C0(n3152), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[224]) );
  XOR2X1 U2201 ( .A(n3153), .B(n3154), .Y(n3152) );
  XOR2X1 U2202 ( .A(n2965), .B(n2983), .Y(n3154) );
  MXI2X1 U2203 ( .A(n3155), .B(n3156), .S0(n375), .Y(n2965) );
  OAI21X1 U2204 ( .A0(n1274), .A1(n1985), .B0(n3157), .Y(n3156) );
  MXI2X1 U2205 ( .A(n3158), .B(n3159), .S0(n2841), .Y(n3157) );
  OAI21X1 U2206 ( .A0(n1985), .A1(n417), .B0(n3160), .Y(n3155) );
  MXI2X1 U2207 ( .A(n3159), .B(n3158), .S0(n2841), .Y(n3160) );
  CLKINVX1 U2208 ( .A(n1987), .Y(n2841) );
  XNOR2X1 U2209 ( .A(n1274), .B(n448), .Y(n1987) );
  NOR2X1 U2210 ( .A(n1465), .B(n1401), .Y(n3158) );
  CLKINVX1 U2211 ( .A(n2839), .Y(n3159) );
  CLKNAND2X2 U2212 ( .A(n1401), .B(n1465), .Y(n2839) );
  CLKINVX1 U2213 ( .A(n3161), .Y(n1985) );
  AOI21X1 U2214 ( .A0(n919), .A1(n1465), .B0(n861), .Y(n3151) );
  AOI21X1 U2215 ( .A0(n1176), .A1(n931), .B0(n959), .Y(n3150) );
  OAI222X1 U2216 ( .A0(n1464), .A1(n3162), .B0(n1051), .B1(n3163), .C0(n3164), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[223]) );
  XOR2X1 U2217 ( .A(n3165), .B(n3166), .Y(n3164) );
  XOR2X1 U2218 ( .A(n2971), .B(n2989), .Y(n3166) );
  MXI2X1 U2219 ( .A(n3167), .B(n3168), .S0(n1528), .Y(n2971) );
  OAI21X1 U2220 ( .A0(n1992), .A1(n418), .B0(n3169), .Y(n3168) );
  MXI2X1 U2221 ( .A(n3170), .B(n3171), .S0(n1994), .Y(n3169) );
  OAI21X1 U2222 ( .A0(n1273), .A1(n1992), .B0(n3172), .Y(n3167) );
  MXI2X1 U2223 ( .A(n3171), .B(n3170), .S0(n1994), .Y(n3172) );
  CLKINVX1 U2224 ( .A(n2959), .Y(n1994) );
  XNOR2X1 U2225 ( .A(n1273), .B(n449), .Y(n2959) );
  CLKINVX1 U2226 ( .A(n2862), .Y(n3170) );
  CLKNAND2X2 U2227 ( .A(n1400), .B(n1464), .Y(n2862) );
  NOR2X1 U2228 ( .A(n1464), .B(n1400), .Y(n3171) );
  CLKINVX1 U2229 ( .A(n3173), .Y(n1992) );
  AOI21X1 U2230 ( .A0(n919), .A1(n1464), .B0(n861), .Y(n3163) );
  AOI21X1 U2231 ( .A0(n1051), .A1(n931), .B0(n959), .Y(n3162) );
  OAI222X1 U2232 ( .A0(n1463), .A1(n3174), .B0(n1055), .B1(n3175), .C0(n3176), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[222]) );
  XOR2X1 U2233 ( .A(n3177), .B(n3178), .Y(n3176) );
  XOR2X1 U2234 ( .A(n2977), .B(n2995), .Y(n3178) );
  MXI2X1 U2235 ( .A(n3179), .B(n3180), .S0(n1527), .Y(n2977) );
  OAI21X1 U2236 ( .A0(n1999), .A1(n419), .B0(n3181), .Y(n3180) );
  MXI2X1 U2237 ( .A(n3182), .B(n3183), .S0(n2001), .Y(n3181) );
  OAI21X1 U2238 ( .A0(n1272), .A1(n1999), .B0(n3184), .Y(n3179) );
  MXI2X1 U2239 ( .A(n3183), .B(n3182), .S0(n2001), .Y(n3184) );
  CLKINVX1 U2240 ( .A(n3023), .Y(n2001) );
  XNOR2X1 U2241 ( .A(n1272), .B(n450), .Y(n3023) );
  CLKINVX1 U2242 ( .A(n2877), .Y(n3182) );
  CLKNAND2X2 U2243 ( .A(n1399), .B(n1463), .Y(n2877) );
  NOR2X1 U2244 ( .A(n1463), .B(n1399), .Y(n3183) );
  CLKINVX1 U2245 ( .A(n3185), .Y(n1999) );
  AOI21X1 U2246 ( .A0(n919), .A1(n1463), .B0(n866), .Y(n3175) );
  AOI21X1 U2247 ( .A0(n1055), .A1(n931), .B0(n959), .Y(n3174) );
  OAI222X1 U2248 ( .A0(n1462), .A1(n3186), .B0(n1059), .B1(n3187), .C0(n3188), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[221]) );
  XNOR2X1 U2249 ( .A(n3189), .B(n3190), .Y(n3188) );
  XOR2X1 U2250 ( .A(n2983), .B(n3001), .Y(n3190) );
  MXI2X1 U2251 ( .A(n3191), .B(n3192), .S0(n1526), .Y(n2983) );
  OAI21X1 U2252 ( .A0(n2006), .A1(n420), .B0(n3193), .Y(n3192) );
  MXI2X1 U2253 ( .A(n3194), .B(n3195), .S0(n2008), .Y(n3193) );
  OAI21X1 U2254 ( .A0(n1271), .A1(n2006), .B0(n3196), .Y(n3191) );
  MXI2X1 U2255 ( .A(n3195), .B(n3194), .S0(n2008), .Y(n3196) );
  CLKINVX1 U2256 ( .A(n3090), .Y(n2008) );
  XNOR2X1 U2257 ( .A(n1271), .B(n451), .Y(n3090) );
  CLKINVX1 U2258 ( .A(n2894), .Y(n3194) );
  CLKNAND2X2 U2259 ( .A(n1398), .B(n1462), .Y(n2894) );
  NOR2X1 U2260 ( .A(n1462), .B(n1398), .Y(n3195) );
  CLKINVX1 U2261 ( .A(n3197), .Y(n2006) );
  AOI21X1 U2262 ( .A0(n919), .A1(n1462), .B0(n861), .Y(n3187) );
  AOI21X1 U2263 ( .A0(n1059), .A1(n931), .B0(n959), .Y(n3186) );
  OAI222X1 U2264 ( .A0(n1461), .A1(n3198), .B0(n1063), .B1(n3199), .C0(n3200), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[220]) );
  XNOR2X1 U2265 ( .A(n3201), .B(n3202), .Y(n3200) );
  XOR2X1 U2266 ( .A(n2989), .B(n3007), .Y(n3202) );
  MXI2X1 U2267 ( .A(n3203), .B(n3204), .S0(n1525), .Y(n2989) );
  OAI21X1 U2268 ( .A0(n2013), .A1(n421), .B0(n3205), .Y(n3204) );
  MXI2X1 U2269 ( .A(n3206), .B(n3207), .S0(n2015), .Y(n3205) );
  OAI21X1 U2270 ( .A0(n1270), .A1(n2013), .B0(n3208), .Y(n3203) );
  MXI2X1 U2271 ( .A(n3207), .B(n3206), .S0(n2015), .Y(n3208) );
  CLKINVX1 U2272 ( .A(n3209), .Y(n2015) );
  CLKINVX1 U2273 ( .A(n2913), .Y(n3206) );
  CLKNAND2X2 U2274 ( .A(n1397), .B(n1461), .Y(n2913) );
  NOR2X1 U2275 ( .A(n1461), .B(n1397), .Y(n3207) );
  CLKINVX1 U2276 ( .A(n3210), .Y(n2013) );
  AOI21X1 U2277 ( .A0(n919), .A1(n1461), .B0(n861), .Y(n3199) );
  AOI21X1 U2278 ( .A0(n1063), .A1(n931), .B0(n959), .Y(n3198) );
  OAI222X1 U2279 ( .A0(n877), .A1(n3211), .B0(n903), .B1(n3212), .C0(n856), 
        .C1(n1720), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[21]) );
  XOR2X1 U2280 ( .A(n2213), .B(n3213), .Y(n3212) );
  XOR2X1 U2281 ( .A(n2181), .B(n2116), .Y(n3213) );
  MXI2X1 U2282 ( .A(n2479), .B(n3214), .S0(n1495), .Y(n2116) );
  XOR2X1 U2283 ( .A(n1367), .B(n354), .Y(n2479) );
  MXI2X1 U2284 ( .A(n2912), .B(n3209), .S0(n1461), .Y(n2181) );
  XNOR2X1 U2285 ( .A(n1270), .B(n452), .Y(n3209) );
  XNOR2X1 U2286 ( .A(n1333), .B(n1525), .Y(n2912) );
  OAI222X1 U2287 ( .A0(n1460), .A1(n3215), .B0(n1067), .B1(n3216), .C0(n3217), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[219]) );
  XNOR2X1 U2288 ( .A(n3218), .B(n3219), .Y(n3217) );
  XOR2X1 U2289 ( .A(n2995), .B(n3013), .Y(n3219) );
  MXI2X1 U2290 ( .A(n3220), .B(n3221), .S0(n1524), .Y(n2995) );
  OAI21X1 U2291 ( .A0(n2020), .A1(n422), .B0(n3222), .Y(n3221) );
  MXI2X1 U2292 ( .A(n3223), .B(n3224), .S0(n2022), .Y(n3222) );
  OAI21X1 U2293 ( .A0(n1269), .A1(n2020), .B0(n3225), .Y(n3220) );
  MXI2X1 U2294 ( .A(n3224), .B(n3223), .S0(n2022), .Y(n3225) );
  CLKINVX1 U2295 ( .A(n3226), .Y(n2022) );
  CLKINVX1 U2296 ( .A(n2767), .Y(n3223) );
  CLKNAND2X2 U2297 ( .A(n1396), .B(n1460), .Y(n2767) );
  NOR2X1 U2298 ( .A(n1460), .B(n1396), .Y(n3224) );
  CLKINVX1 U2299 ( .A(n3227), .Y(n2020) );
  AOI21X1 U2300 ( .A0(n919), .A1(n1460), .B0(n862), .Y(n3216) );
  AOI21X1 U2301 ( .A0(n1067), .A1(n931), .B0(n959), .Y(n3215) );
  OAI222X1 U2302 ( .A0(n1459), .A1(n3228), .B0(n1071), .B1(n3229), .C0(n3230), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[218]) );
  XNOR2X1 U2303 ( .A(n3231), .B(n3232), .Y(n3230) );
  XOR2X1 U2304 ( .A(n3001), .B(n3019), .Y(n3232) );
  MXI2X1 U2305 ( .A(n3233), .B(n3234), .S0(n1523), .Y(n3001) );
  OAI21X1 U2306 ( .A0(n2027), .A1(n423), .B0(n3235), .Y(n3234) );
  MXI2X1 U2307 ( .A(n3236), .B(n3237), .S0(n2029), .Y(n3235) );
  OAI21X1 U2308 ( .A0(n1268), .A1(n2027), .B0(n3238), .Y(n3233) );
  MXI2X1 U2309 ( .A(n3237), .B(n3236), .S0(n2029), .Y(n3238) );
  CLKINVX1 U2310 ( .A(n3239), .Y(n2029) );
  CLKINVX1 U2311 ( .A(n2787), .Y(n3236) );
  CLKNAND2X2 U2312 ( .A(n1395), .B(n1459), .Y(n2787) );
  NOR2X1 U2313 ( .A(n1459), .B(n1395), .Y(n3237) );
  CLKINVX1 U2314 ( .A(n3240), .Y(n2027) );
  AOI21X1 U2315 ( .A0(n920), .A1(n1459), .B0(n862), .Y(n3229) );
  AOI21X1 U2316 ( .A0(n1071), .A1(n932), .B0(n958), .Y(n3228) );
  OAI222X1 U2317 ( .A0(n1458), .A1(n3241), .B0(n1075), .B1(n3242), .C0(n3243), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[217]) );
  XNOR2X1 U2318 ( .A(n3244), .B(n3245), .Y(n3243) );
  XOR2X1 U2319 ( .A(n3007), .B(n3029), .Y(n3245) );
  MXI2X1 U2320 ( .A(n3246), .B(n3247), .S0(n1522), .Y(n3007) );
  OAI21X1 U2321 ( .A0(n2034), .A1(n424), .B0(n3248), .Y(n3247) );
  MXI2X1 U2322 ( .A(n3249), .B(n3250), .S0(n2036), .Y(n3248) );
  OAI21X1 U2323 ( .A0(n1267), .A1(n2034), .B0(n3251), .Y(n3246) );
  MXI2X1 U2324 ( .A(n3250), .B(n3249), .S0(n2036), .Y(n3251) );
  CLKINVX1 U2325 ( .A(n3252), .Y(n2036) );
  CLKINVX1 U2326 ( .A(n2803), .Y(n3249) );
  CLKNAND2X2 U2327 ( .A(n1394), .B(n1458), .Y(n2803) );
  NOR2X1 U2328 ( .A(n1458), .B(n1394), .Y(n3250) );
  CLKINVX1 U2329 ( .A(n3253), .Y(n2034) );
  AOI21X1 U2330 ( .A0(n920), .A1(n1458), .B0(n862), .Y(n3242) );
  AOI21X1 U2331 ( .A0(n1075), .A1(n932), .B0(n958), .Y(n3241) );
  OAI222X1 U2332 ( .A0(n1457), .A1(n3254), .B0(n1079), .B1(n3255), .C0(n3256), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[216]) );
  XOR2X1 U2333 ( .A(n3035), .B(n3257), .Y(n3256) );
  XOR2X1 U2334 ( .A(n2921), .B(n3013), .Y(n3257) );
  MXI2X1 U2335 ( .A(n3258), .B(n3259), .S0(n1521), .Y(n3013) );
  OAI21X1 U2336 ( .A0(n2041), .A1(n425), .B0(n3260), .Y(n3259) );
  MXI2X1 U2337 ( .A(n3261), .B(n3262), .S0(n2043), .Y(n3260) );
  OAI21X1 U2338 ( .A0(n1266), .A1(n2041), .B0(n3263), .Y(n3258) );
  MXI2X1 U2339 ( .A(n3262), .B(n3261), .S0(n2043), .Y(n3263) );
  CLKINVX1 U2340 ( .A(n3264), .Y(n2043) );
  CLKINVX1 U2341 ( .A(n2819), .Y(n3261) );
  CLKNAND2X2 U2342 ( .A(n1393), .B(n1457), .Y(n2819) );
  NOR2X1 U2343 ( .A(n1457), .B(n1393), .Y(n3262) );
  CLKINVX1 U2344 ( .A(n3265), .Y(n2041) );
  AOI21X1 U2345 ( .A0(n920), .A1(n1457), .B0(n862), .Y(n3255) );
  AOI21X1 U2346 ( .A0(n1079), .A1(n932), .B0(n958), .Y(n3254) );
  OAI222X1 U2347 ( .A0(n1456), .A1(n3266), .B0(n1083), .B1(n3267), .C0(n3268), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[215]) );
  XOR2X1 U2348 ( .A(n3041), .B(n3269), .Y(n3268) );
  XOR2X1 U2349 ( .A(n2929), .B(n3019), .Y(n3269) );
  MXI2X1 U2350 ( .A(n3270), .B(n3271), .S0(n1520), .Y(n3019) );
  OAI21X1 U2351 ( .A0(n2049), .A1(n426), .B0(n3272), .Y(n3271) );
  MXI2X1 U2352 ( .A(n3273), .B(n3274), .S0(n2051), .Y(n3272) );
  OAI21X1 U2353 ( .A0(n1265), .A1(n2049), .B0(n3275), .Y(n3270) );
  MXI2X1 U2354 ( .A(n3274), .B(n3273), .S0(n2051), .Y(n3275) );
  CLKINVX1 U2355 ( .A(n3276), .Y(n2051) );
  CLKINVX1 U2356 ( .A(n2835), .Y(n3273) );
  CLKNAND2X2 U2357 ( .A(n1392), .B(n1456), .Y(n2835) );
  NOR2X1 U2358 ( .A(n1456), .B(n1392), .Y(n3274) );
  CLKINVX1 U2359 ( .A(n3277), .Y(n2049) );
  AOI21X1 U2360 ( .A0(n920), .A1(n1456), .B0(n862), .Y(n3267) );
  AOI21X1 U2361 ( .A0(n1083), .A1(n932), .B0(n958), .Y(n3266) );
  OAI222X1 U2362 ( .A0(n1455), .A1(n3278), .B0(n1087), .B1(n3279), .C0(n3280), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[214]) );
  XOR2X1 U2363 ( .A(n3047), .B(n3281), .Y(n3280) );
  XOR2X1 U2364 ( .A(n2936), .B(n3029), .Y(n3281) );
  MXI2X1 U2365 ( .A(n3282), .B(n3283), .S0(n1519), .Y(n3029) );
  OAI21X1 U2366 ( .A0(n2063), .A1(n427), .B0(n3284), .Y(n3283) );
  MXI2X1 U2367 ( .A(n3285), .B(n3286), .S0(n2065), .Y(n3284) );
  OAI21X1 U2368 ( .A0(n1264), .A1(n2063), .B0(n3287), .Y(n3282) );
  MXI2X1 U2369 ( .A(n3286), .B(n3285), .S0(n2065), .Y(n3287) );
  CLKINVX1 U2370 ( .A(n3288), .Y(n2065) );
  CLKINVX1 U2371 ( .A(n2858), .Y(n3285) );
  CLKNAND2X2 U2372 ( .A(n1391), .B(n1455), .Y(n2858) );
  NOR2X1 U2373 ( .A(n1455), .B(n1391), .Y(n3286) );
  CLKINVX1 U2374 ( .A(n3289), .Y(n2063) );
  AOI21X1 U2375 ( .A0(n920), .A1(n1455), .B0(n862), .Y(n3279) );
  AOI21X1 U2376 ( .A0(n1087), .A1(n932), .B0(n958), .Y(n3278) );
  OAI222X1 U2377 ( .A0(n1454), .A1(n3290), .B0(n1091), .B1(n3291), .C0(n3292), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[213]) );
  XOR2X1 U2378 ( .A(n3053), .B(n3293), .Y(n3292) );
  XOR2X1 U2379 ( .A(n2922), .B(n3035), .Y(n3293) );
  MXI2X1 U2380 ( .A(n3294), .B(n3295), .S0(n1518), .Y(n3035) );
  OAI21X1 U2381 ( .A0(n2071), .A1(n428), .B0(n3296), .Y(n3295) );
  MXI2X1 U2382 ( .A(n3297), .B(n3298), .S0(n2073), .Y(n3296) );
  OAI21X1 U2383 ( .A0(n1263), .A1(n2071), .B0(n3299), .Y(n3294) );
  MXI2X1 U2384 ( .A(n3298), .B(n3297), .S0(n2073), .Y(n3299) );
  CLKINVX1 U2385 ( .A(n3300), .Y(n2073) );
  CLKINVX1 U2386 ( .A(n2873), .Y(n3297) );
  CLKNAND2X2 U2387 ( .A(n1390), .B(n1454), .Y(n2873) );
  NOR2X1 U2388 ( .A(n1454), .B(n1390), .Y(n3298) );
  CLKINVX1 U2389 ( .A(n3301), .Y(n2071) );
  MXI2X1 U2390 ( .A(n3302), .B(n3303), .S0(n358), .Y(n2922) );
  OAI21X1 U2391 ( .A0(n1302), .A1(n3304), .B0(n3305), .Y(n3303) );
  MXI2X1 U2392 ( .A(n3306), .B(n3307), .S0(n2511), .Y(n3305) );
  OAI21X1 U2393 ( .A0(n3304), .A1(n384), .B0(n3308), .Y(n3302) );
  MXI2X1 U2394 ( .A(n3307), .B(n3306), .S0(n2511), .Y(n3308) );
  CLKINVX1 U2395 ( .A(n3309), .Y(n2511) );
  NOR2X1 U2396 ( .A(n1493), .B(n1429), .Y(n3306) );
  CLKINVX1 U2397 ( .A(n2509), .Y(n3307) );
  CLKNAND2X2 U2398 ( .A(n1429), .B(n1493), .Y(n2509) );
  AOI21X1 U2399 ( .A0(n920), .A1(n1454), .B0(n862), .Y(n3291) );
  AOI21X1 U2400 ( .A0(n1091), .A1(n932), .B0(n958), .Y(n3290) );
  OAI222X1 U2401 ( .A0(n1453), .A1(n3310), .B0(n1095), .B1(n3311), .C0(n3312), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[212]) );
  XOR2X1 U2402 ( .A(n3059), .B(n3313), .Y(n3312) );
  XOR2X1 U2403 ( .A(n2930), .B(n3041), .Y(n3313) );
  MXI2X1 U2404 ( .A(n3314), .B(n3315), .S0(n1517), .Y(n3041) );
  OAI21X1 U2405 ( .A0(n2079), .A1(n339), .B0(n3316), .Y(n3315) );
  MXI2X1 U2406 ( .A(n2890), .B(n3317), .S0(n2081), .Y(n3316) );
  OAI21X1 U2407 ( .A0(n1262), .A1(n2079), .B0(n3318), .Y(n3314) );
  MXI2X1 U2408 ( .A(n3317), .B(n2890), .S0(n2081), .Y(n3318) );
  AND2X1 U2409 ( .A(n1389), .B(n1453), .Y(n2890) );
  NOR2X1 U2410 ( .A(n1453), .B(n1389), .Y(n3317) );
  CLKINVX1 U2411 ( .A(n3319), .Y(n2079) );
  MXI2X1 U2412 ( .A(n3320), .B(n3321), .S0(n360), .Y(n2930) );
  OAI21X1 U2413 ( .A0(n1301), .A1(n3322), .B0(n3323), .Y(n3321) );
  MXI2X1 U2414 ( .A(n3324), .B(n3325), .S0(n2522), .Y(n3323) );
  OAI21X1 U2415 ( .A0(n3322), .A1(n385), .B0(n3326), .Y(n3320) );
  MXI2X1 U2416 ( .A(n3325), .B(n3324), .S0(n2522), .Y(n3326) );
  CLKINVX1 U2417 ( .A(n3327), .Y(n2522) );
  NOR2X1 U2418 ( .A(n1492), .B(n1428), .Y(n3324) );
  CLKINVX1 U2419 ( .A(n2520), .Y(n3325) );
  CLKNAND2X2 U2420 ( .A(n1428), .B(n1492), .Y(n2520) );
  AOI21X1 U2421 ( .A0(n920), .A1(n1453), .B0(n863), .Y(n3311) );
  AOI21X1 U2422 ( .A0(n1095), .A1(n932), .B0(n958), .Y(n3310) );
  OAI222X1 U2423 ( .A0(n1452), .A1(n3328), .B0(n1099), .B1(n3329), .C0(n3330), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[211]) );
  XOR2X1 U2424 ( .A(n3063), .B(n3331), .Y(n3330) );
  XOR2X1 U2425 ( .A(n2937), .B(n3047), .Y(n3331) );
  MXI2X1 U2426 ( .A(n3332), .B(n3333), .S0(n1516), .Y(n3047) );
  OAI21X1 U2427 ( .A0(n2087), .A1(n340), .B0(n3334), .Y(n3333) );
  MXI2X1 U2428 ( .A(n2909), .B(n3335), .S0(n2089), .Y(n3334) );
  OAI21X1 U2429 ( .A0(n1261), .A1(n2087), .B0(n3336), .Y(n3332) );
  MXI2X1 U2430 ( .A(n3335), .B(n2909), .S0(n2089), .Y(n3336) );
  AND2X1 U2431 ( .A(n1388), .B(n1452), .Y(n2909) );
  NOR2X1 U2432 ( .A(n1452), .B(n1388), .Y(n3335) );
  CLKINVX1 U2433 ( .A(n3337), .Y(n2087) );
  MXI2X1 U2434 ( .A(n3338), .B(n3339), .S0(n362), .Y(n2937) );
  OAI21X1 U2435 ( .A0(n1300), .A1(n3340), .B0(n3341), .Y(n3339) );
  MXI2X1 U2436 ( .A(n3342), .B(n3343), .S0(n2531), .Y(n3341) );
  OAI21X1 U2437 ( .A0(n3340), .A1(n386), .B0(n3344), .Y(n3338) );
  MXI2X1 U2438 ( .A(n3343), .B(n3342), .S0(n2531), .Y(n3344) );
  CLKINVX1 U2439 ( .A(n3345), .Y(n2531) );
  NOR2X1 U2440 ( .A(n1491), .B(n1427), .Y(n3342) );
  CLKINVX1 U2441 ( .A(n2529), .Y(n3343) );
  CLKNAND2X2 U2442 ( .A(n1427), .B(n1491), .Y(n2529) );
  AOI21X1 U2443 ( .A0(n920), .A1(n1452), .B0(n863), .Y(n3329) );
  AOI21X1 U2444 ( .A0(n1099), .A1(n932), .B0(n958), .Y(n3328) );
  OAI222X1 U2445 ( .A0(n1451), .A1(n3346), .B0(n1103), .B1(n3347), .C0(n3348), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[210]) );
  XOR2X1 U2446 ( .A(n3068), .B(n3349), .Y(n3348) );
  XOR2X1 U2447 ( .A(n2941), .B(n3053), .Y(n3349) );
  MXI2X1 U2448 ( .A(n3350), .B(n3351), .S0(n1515), .Y(n3053) );
  OAI21X1 U2449 ( .A0(n2095), .A1(n429), .B0(n3352), .Y(n3351) );
  MXI2X1 U2450 ( .A(n3353), .B(n3354), .S0(n2097), .Y(n3352) );
  OAI21X1 U2451 ( .A0(n1260), .A1(n2095), .B0(n3355), .Y(n3350) );
  MXI2X1 U2452 ( .A(n3354), .B(n3353), .S0(n2097), .Y(n3355) );
  CLKINVX1 U2453 ( .A(n3356), .Y(n2097) );
  CLKINVX1 U2454 ( .A(n2640), .Y(n3353) );
  CLKNAND2X2 U2455 ( .A(n1387), .B(n1451), .Y(n2640) );
  NOR2X1 U2456 ( .A(n1451), .B(n1387), .Y(n3354) );
  CLKINVX1 U2457 ( .A(n3357), .Y(n2095) );
  MXI2X1 U2458 ( .A(n3358), .B(n3359), .S0(n344), .Y(n2941) );
  OAI21X1 U2459 ( .A0(n1299), .A1(n3360), .B0(n3361), .Y(n3359) );
  MXI2X1 U2460 ( .A(n3362), .B(n3363), .S0(n2540), .Y(n3361) );
  OAI21X1 U2461 ( .A0(n3360), .A1(n387), .B0(n3364), .Y(n3358) );
  MXI2X1 U2462 ( .A(n3363), .B(n3362), .S0(n2540), .Y(n3364) );
  CLKINVX1 U2463 ( .A(n3365), .Y(n2540) );
  NOR2X1 U2464 ( .A(n1490), .B(n1426), .Y(n3362) );
  CLKINVX1 U2465 ( .A(n2538), .Y(n3363) );
  CLKNAND2X2 U2466 ( .A(n1426), .B(n1490), .Y(n2538) );
  AOI21X1 U2467 ( .A0(n920), .A1(n1451), .B0(n863), .Y(n3347) );
  AOI21X1 U2468 ( .A0(n1103), .A1(n933), .B0(n958), .Y(n3346) );
  OAI222X1 U2469 ( .A0(n877), .A1(n3366), .B0(n902), .B1(n3367), .C0(n856), 
        .C1(n1719), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[20]) );
  XNOR2X1 U2470 ( .A(n2219), .B(n3368), .Y(n3367) );
  XOR2X1 U2471 ( .A(n2184), .B(n2122), .Y(n3368) );
  MXI2X1 U2472 ( .A(n2498), .B(n3369), .S0(n1494), .Y(n2122) );
  XOR2X1 U2473 ( .A(n1366), .B(n356), .Y(n2498) );
  MXI2X1 U2474 ( .A(n2766), .B(n3226), .S0(n1460), .Y(n2184) );
  XNOR2X1 U2475 ( .A(n1269), .B(n453), .Y(n3226) );
  XNOR2X1 U2476 ( .A(n1332), .B(n1524), .Y(n2766) );
  OAI222X1 U2477 ( .A0(n1450), .A1(n3370), .B0(n1107), .B1(n3371), .C0(n3372), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[209]) );
  XOR2X1 U2478 ( .A(n3073), .B(n3373), .Y(n3372) );
  XOR2X1 U2479 ( .A(n2947), .B(n3059), .Y(n3373) );
  MXI2X1 U2480 ( .A(n3374), .B(n3375), .S0(n1514), .Y(n3059) );
  OAI21X1 U2481 ( .A0(n2103), .A1(n430), .B0(n3376), .Y(n3375) );
  MXI2X1 U2482 ( .A(n3377), .B(n3378), .S0(n2105), .Y(n3376) );
  OAI21X1 U2483 ( .A0(n1259), .A1(n2103), .B0(n3379), .Y(n3374) );
  MXI2X1 U2484 ( .A(n3378), .B(n3377), .S0(n2105), .Y(n3379) );
  CLKINVX1 U2485 ( .A(n3380), .Y(n2105) );
  CLKINVX1 U2486 ( .A(n2651), .Y(n3377) );
  CLKNAND2X2 U2487 ( .A(n1386), .B(n1450), .Y(n2651) );
  NOR2X1 U2488 ( .A(n1450), .B(n1386), .Y(n3378) );
  CLKINVX1 U2489 ( .A(n3381), .Y(n2103) );
  MXI2X1 U2490 ( .A(n3382), .B(n3383), .S0(n345), .Y(n2947) );
  OAI21X1 U2491 ( .A0(n1298), .A1(n3384), .B0(n3385), .Y(n3383) );
  MXI2X1 U2492 ( .A(n3386), .B(n3387), .S0(n2549), .Y(n3385) );
  OAI21X1 U2493 ( .A0(n3384), .A1(n388), .B0(n3388), .Y(n3382) );
  MXI2X1 U2494 ( .A(n3387), .B(n3386), .S0(n2549), .Y(n3388) );
  CLKINVX1 U2495 ( .A(n3389), .Y(n2549) );
  NOR2X1 U2496 ( .A(n1489), .B(n1425), .Y(n3386) );
  CLKINVX1 U2497 ( .A(n2547), .Y(n3387) );
  CLKNAND2X2 U2498 ( .A(n1425), .B(n1489), .Y(n2547) );
  AOI21X1 U2499 ( .A0(n920), .A1(n1450), .B0(n863), .Y(n3371) );
  AOI21X1 U2500 ( .A0(n1107), .A1(n933), .B0(n958), .Y(n3370) );
  OAI222X1 U2501 ( .A0(n1449), .A1(n3390), .B0(n1111), .B1(n3391), .C0(n3392), 
        .C1(n895), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[208]) );
  XOR2X1 U2502 ( .A(n3078), .B(n3393), .Y(n3392) );
  XOR2X1 U2503 ( .A(n2953), .B(n3063), .Y(n3393) );
  MXI2X1 U2504 ( .A(n3394), .B(n3395), .S0(n348), .Y(n3063) );
  OAI21X1 U2505 ( .A0(n1258), .A1(n3396), .B0(n3397), .Y(n3395) );
  MXI2X1 U2506 ( .A(n3398), .B(n3399), .S0(n2664), .Y(n3397) );
  OAI21X1 U2507 ( .A0(n3396), .A1(n406), .B0(n3400), .Y(n3394) );
  MXI2X1 U2508 ( .A(n3399), .B(n3398), .S0(n2664), .Y(n3400) );
  CLKINVX1 U2509 ( .A(n3401), .Y(n2664) );
  NOR2X1 U2510 ( .A(n1449), .B(n1385), .Y(n3398) );
  CLKINVX1 U2511 ( .A(n2662), .Y(n3399) );
  CLKNAND2X2 U2512 ( .A(n1385), .B(n1449), .Y(n2662) );
  MXI2X1 U2513 ( .A(n3402), .B(n3403), .S0(n346), .Y(n2953) );
  OAI21X1 U2514 ( .A0(n1297), .A1(n3404), .B0(n3405), .Y(n3403) );
  MXI2X1 U2515 ( .A(n3406), .B(n3407), .S0(n2557), .Y(n3405) );
  OAI21X1 U2516 ( .A0(n3404), .A1(n389), .B0(n3408), .Y(n3402) );
  MXI2X1 U2517 ( .A(n3407), .B(n3406), .S0(n2557), .Y(n3408) );
  CLKINVX1 U2518 ( .A(n3409), .Y(n2557) );
  NOR2X1 U2519 ( .A(n1488), .B(n1424), .Y(n3406) );
  CLKINVX1 U2520 ( .A(n2555), .Y(n3407) );
  CLKNAND2X2 U2521 ( .A(n1424), .B(n1488), .Y(n2555) );
  AOI21X1 U2522 ( .A0(n920), .A1(n1449), .B0(n863), .Y(n3391) );
  AOI21X1 U2523 ( .A0(n1111), .A1(n933), .B0(n958), .Y(n3390) );
  OAI222X1 U2524 ( .A0(n1448), .A1(n3410), .B0(n1115), .B1(n3411), .C0(n3412), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[207]) );
  XOR2X1 U2525 ( .A(n3094), .B(n3413), .Y(n3412) );
  XOR2X1 U2526 ( .A(n2963), .B(n3068), .Y(n3413) );
  MXI2X1 U2527 ( .A(n3414), .B(n3415), .S0(n349), .Y(n3068) );
  OAI21X1 U2528 ( .A0(n1257), .A1(n3416), .B0(n3417), .Y(n3415) );
  MXI2X1 U2529 ( .A(n3418), .B(n3419), .S0(n2679), .Y(n3417) );
  OAI21X1 U2530 ( .A0(n3416), .A1(n407), .B0(n3420), .Y(n3414) );
  MXI2X1 U2531 ( .A(n3419), .B(n3418), .S0(n2679), .Y(n3420) );
  CLKINVX1 U2532 ( .A(n3421), .Y(n2679) );
  NOR2X1 U2533 ( .A(n1448), .B(n1384), .Y(n3418) );
  CLKINVX1 U2534 ( .A(n2677), .Y(n3419) );
  CLKNAND2X2 U2535 ( .A(n1384), .B(n1448), .Y(n2677) );
  MXI2X1 U2536 ( .A(n3422), .B(n3423), .S0(n1551), .Y(n2963) );
  OAI21X1 U2537 ( .A0(n3424), .A1(n390), .B0(n3425), .Y(n3423) );
  MXI2X1 U2538 ( .A(n3426), .B(n3427), .S0(n2565), .Y(n3425) );
  OAI21X1 U2539 ( .A0(n1296), .A1(n3424), .B0(n3428), .Y(n3422) );
  MXI2X1 U2540 ( .A(n3427), .B(n3426), .S0(n2565), .Y(n3428) );
  CLKINVX1 U2541 ( .A(n3429), .Y(n2565) );
  CLKINVX1 U2542 ( .A(n2563), .Y(n3426) );
  CLKNAND2X2 U2543 ( .A(n1423), .B(n1487), .Y(n2563) );
  NOR2X1 U2544 ( .A(n1487), .B(n1423), .Y(n3427) );
  AOI21X1 U2545 ( .A0(n920), .A1(n1448), .B0(n863), .Y(n3411) );
  AOI21X1 U2546 ( .A0(n1115), .A1(n933), .B0(n958), .Y(n3410) );
  OAI222X1 U2547 ( .A0(n1447), .A1(n3430), .B0(n1119), .B1(n3431), .C0(n3432), 
        .C1(n894), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[206]) );
  XOR2X1 U2548 ( .A(n3105), .B(n3433), .Y(n3432) );
  XOR2X1 U2549 ( .A(n2969), .B(n3073), .Y(n3433) );
  MXI2X1 U2550 ( .A(n3434), .B(n3435), .S0(n371), .Y(n3073) );
  OAI21X1 U2551 ( .A0(n1256), .A1(n3436), .B0(n3437), .Y(n3435) );
  MXI2X1 U2552 ( .A(n3438), .B(n3439), .S0(n2692), .Y(n3437) );
  OAI21X1 U2553 ( .A0(n3436), .A1(n408), .B0(n3440), .Y(n3434) );
  MXI2X1 U2554 ( .A(n3439), .B(n3438), .S0(n2692), .Y(n3440) );
  CLKINVX1 U2555 ( .A(n3441), .Y(n2692) );
  NOR2X1 U2556 ( .A(n1447), .B(n1383), .Y(n3438) );
  CLKINVX1 U2557 ( .A(n2690), .Y(n3439) );
  CLKNAND2X2 U2558 ( .A(n1383), .B(n1447), .Y(n2690) );
  MXI2X1 U2559 ( .A(n3442), .B(n3443), .S0(n347), .Y(n2969) );
  OAI21X1 U2560 ( .A0(n1295), .A1(n3444), .B0(n3445), .Y(n3443) );
  MXI2X1 U2561 ( .A(n3446), .B(n3447), .S0(n2573), .Y(n3445) );
  OAI21X1 U2562 ( .A0(n3444), .A1(n391), .B0(n3448), .Y(n3442) );
  MXI2X1 U2563 ( .A(n3447), .B(n3446), .S0(n2573), .Y(n3448) );
  CLKINVX1 U2564 ( .A(n3449), .Y(n2573) );
  NOR2X1 U2565 ( .A(n1486), .B(n1422), .Y(n3446) );
  CLKINVX1 U2566 ( .A(n2571), .Y(n3447) );
  CLKNAND2X2 U2567 ( .A(n1422), .B(n1486), .Y(n2571) );
  AOI21X1 U2568 ( .A0(n921), .A1(n1447), .B0(n863), .Y(n3431) );
  AOI21X1 U2569 ( .A0(n1119), .A1(n933), .B0(n958), .Y(n3430) );
  OAI222X1 U2570 ( .A0(n1446), .A1(n3450), .B0(n1123), .B1(n3451), .C0(n3452), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[205]) );
  XOR2X1 U2571 ( .A(n3117), .B(n3453), .Y(n3452) );
  XOR2X1 U2572 ( .A(n2975), .B(n3078), .Y(n3453) );
  MXI2X1 U2573 ( .A(n3454), .B(n3455), .S0(n1510), .Y(n3078) );
  OAI21X1 U2574 ( .A0(n3456), .A1(n431), .B0(n3457), .Y(n3455) );
  MXI2X1 U2575 ( .A(n3458), .B(n3459), .S0(n2712), .Y(n3457) );
  OAI21X1 U2576 ( .A0(n1255), .A1(n3456), .B0(n3460), .Y(n3454) );
  MXI2X1 U2577 ( .A(n3459), .B(n3458), .S0(n2712), .Y(n3460) );
  CLKINVX1 U2578 ( .A(n2710), .Y(n3458) );
  CLKNAND2X2 U2579 ( .A(n1382), .B(n1446), .Y(n2710) );
  NOR2X1 U2580 ( .A(n1446), .B(n1382), .Y(n3459) );
  MXI2X1 U2581 ( .A(n3461), .B(n3462), .S0(n359), .Y(n2975) );
  OAI21X1 U2582 ( .A0(n1294), .A1(n3463), .B0(n3464), .Y(n3462) );
  MXI2X1 U2583 ( .A(n3465), .B(n3466), .S0(n2583), .Y(n3464) );
  OAI21X1 U2584 ( .A0(n3463), .A1(n392), .B0(n3467), .Y(n3461) );
  MXI2X1 U2585 ( .A(n3466), .B(n3465), .S0(n2583), .Y(n3467) );
  CLKINVX1 U2586 ( .A(n3468), .Y(n2583) );
  NOR2X1 U2587 ( .A(n1485), .B(n1421), .Y(n3465) );
  CLKINVX1 U2588 ( .A(n2581), .Y(n3466) );
  CLKNAND2X2 U2589 ( .A(n1421), .B(n1485), .Y(n2581) );
  AOI21X1 U2590 ( .A0(n921), .A1(n1446), .B0(n864), .Y(n3451) );
  AOI21X1 U2591 ( .A0(n1123), .A1(n933), .B0(n957), .Y(n3450) );
  OAI222X1 U2592 ( .A0(n1445), .A1(n3469), .B0(n1127), .B1(n3470), .C0(n3471), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[204]) );
  XOR2X1 U2593 ( .A(n3129), .B(n3472), .Y(n3471) );
  XOR2X1 U2594 ( .A(n2981), .B(n3094), .Y(n3472) );
  MXI2X1 U2595 ( .A(n3473), .B(n3474), .S0(n1509), .Y(n3094) );
  OAI21X1 U2596 ( .A0(n3475), .A1(n432), .B0(n3476), .Y(n3474) );
  MXI2X1 U2597 ( .A(n3477), .B(n3478), .S0(n2724), .Y(n3476) );
  OAI21X1 U2598 ( .A0(n1254), .A1(n3475), .B0(n3479), .Y(n3473) );
  MXI2X1 U2599 ( .A(n3478), .B(n3477), .S0(n2724), .Y(n3479) );
  CLKINVX1 U2600 ( .A(n2722), .Y(n3477) );
  CLKNAND2X2 U2601 ( .A(n1381), .B(n1445), .Y(n2722) );
  NOR2X1 U2602 ( .A(n1445), .B(n1381), .Y(n3478) );
  MXI2X1 U2603 ( .A(n3480), .B(n3481), .S0(n361), .Y(n2981) );
  OAI21X1 U2604 ( .A0(n1293), .A1(n3482), .B0(n3483), .Y(n3481) );
  MXI2X1 U2605 ( .A(n3484), .B(n3485), .S0(n2602), .Y(n3483) );
  OAI21X1 U2606 ( .A0(n3482), .A1(n393), .B0(n3486), .Y(n3480) );
  MXI2X1 U2607 ( .A(n3485), .B(n3484), .S0(n2602), .Y(n3486) );
  CLKINVX1 U2608 ( .A(n3487), .Y(n2602) );
  NOR2X1 U2609 ( .A(n1484), .B(n1420), .Y(n3484) );
  CLKINVX1 U2610 ( .A(n2600), .Y(n3485) );
  CLKNAND2X2 U2611 ( .A(n1420), .B(n1484), .Y(n2600) );
  AOI21X1 U2612 ( .A0(n921), .A1(n1445), .B0(n864), .Y(n3470) );
  AOI21X1 U2613 ( .A0(n1127), .A1(n933), .B0(n957), .Y(n3469) );
  OAI222X1 U2614 ( .A0(n1444), .A1(n3488), .B0(n1131), .B1(n3489), .C0(n3490), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[203]) );
  XOR2X1 U2615 ( .A(n3141), .B(n3491), .Y(n3490) );
  XOR2X1 U2616 ( .A(n2987), .B(n3105), .Y(n3491) );
  MXI2X1 U2617 ( .A(n3492), .B(n3493), .S0(n1508), .Y(n3105) );
  OAI21X1 U2618 ( .A0(n3494), .A1(n433), .B0(n3495), .Y(n3493) );
  MXI2X1 U2619 ( .A(n3496), .B(n3497), .S0(n2735), .Y(n3495) );
  OAI21X1 U2620 ( .A0(n1253), .A1(n3494), .B0(n3498), .Y(n3492) );
  MXI2X1 U2621 ( .A(n3497), .B(n3496), .S0(n2735), .Y(n3498) );
  CLKINVX1 U2622 ( .A(n2733), .Y(n3496) );
  CLKNAND2X2 U2623 ( .A(n1380), .B(n1444), .Y(n2733) );
  NOR2X1 U2624 ( .A(n1444), .B(n1380), .Y(n3497) );
  MXI2X1 U2625 ( .A(n3499), .B(n3500), .S0(n364), .Y(n2987) );
  OAI21X1 U2626 ( .A0(n1292), .A1(n3501), .B0(n3502), .Y(n3500) );
  MXI2X1 U2627 ( .A(n3503), .B(n3504), .S0(n2609), .Y(n3502) );
  OAI21X1 U2628 ( .A0(n3501), .A1(n394), .B0(n3505), .Y(n3499) );
  MXI2X1 U2629 ( .A(n3504), .B(n3503), .S0(n2609), .Y(n3505) );
  CLKINVX1 U2630 ( .A(n2222), .Y(n2609) );
  NOR2X1 U2631 ( .A(n1483), .B(n1419), .Y(n3503) );
  CLKINVX1 U2632 ( .A(n2607), .Y(n3504) );
  CLKNAND2X2 U2633 ( .A(n1419), .B(n1483), .Y(n2607) );
  AOI21X1 U2634 ( .A0(n921), .A1(n1444), .B0(n864), .Y(n3489) );
  AOI21X1 U2635 ( .A0(n1131), .A1(n933), .B0(n957), .Y(n3488) );
  OAI222X1 U2636 ( .A0(n1443), .A1(n3506), .B0(n1135), .B1(n3507), .C0(n3508), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[202]) );
  XOR2X1 U2637 ( .A(n3153), .B(n3509), .Y(n3508) );
  XOR2X1 U2638 ( .A(n2993), .B(n3117), .Y(n3509) );
  MXI2X1 U2639 ( .A(n3510), .B(n3511), .S0(n1507), .Y(n3117) );
  OAI21X1 U2640 ( .A0(n3512), .A1(n434), .B0(n3513), .Y(n3511) );
  MXI2X1 U2641 ( .A(n3514), .B(n3515), .S0(n2746), .Y(n3513) );
  OAI21X1 U2642 ( .A0(n1252), .A1(n3512), .B0(n3516), .Y(n3510) );
  MXI2X1 U2643 ( .A(n3515), .B(n3514), .S0(n2746), .Y(n3516) );
  CLKINVX1 U2644 ( .A(n2744), .Y(n3514) );
  CLKNAND2X2 U2645 ( .A(n1379), .B(n1443), .Y(n2744) );
  NOR2X1 U2646 ( .A(n1443), .B(n1379), .Y(n3515) );
  MXI2X1 U2647 ( .A(n3517), .B(n3518), .S0(n365), .Y(n2993) );
  OAI21X1 U2648 ( .A0(n1291), .A1(n3519), .B0(n3520), .Y(n3518) );
  MXI2X1 U2649 ( .A(n3521), .B(n3522), .S0(n2616), .Y(n3520) );
  OAI21X1 U2650 ( .A0(n3519), .A1(n395), .B0(n3523), .Y(n3517) );
  MXI2X1 U2651 ( .A(n3522), .B(n3521), .S0(n2616), .Y(n3523) );
  CLKINVX1 U2652 ( .A(n2229), .Y(n2616) );
  NOR2X1 U2653 ( .A(n1482), .B(n1418), .Y(n3521) );
  CLKINVX1 U2654 ( .A(n2614), .Y(n3522) );
  CLKNAND2X2 U2655 ( .A(n1418), .B(n1482), .Y(n2614) );
  AOI21X1 U2656 ( .A0(n921), .A1(n1443), .B0(n864), .Y(n3507) );
  AOI21X1 U2657 ( .A0(n1135), .A1(n933), .B0(n957), .Y(n3506) );
  OAI222X1 U2658 ( .A0(n1442), .A1(n3524), .B0(n1139), .B1(n3525), .C0(n3526), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[201]) );
  XOR2X1 U2659 ( .A(n3165), .B(n3527), .Y(n3526) );
  XOR2X1 U2660 ( .A(n2999), .B(n3129), .Y(n3527) );
  MXI2X1 U2661 ( .A(n3528), .B(n3529), .S0(n372), .Y(n3129) );
  OAI21X1 U2662 ( .A0(n1251), .A1(n3530), .B0(n3531), .Y(n3529) );
  MXI2X1 U2663 ( .A(n3532), .B(n3533), .S0(n2756), .Y(n3531) );
  OAI21X1 U2664 ( .A0(n3530), .A1(n409), .B0(n3534), .Y(n3528) );
  MXI2X1 U2665 ( .A(n3533), .B(n3532), .S0(n2756), .Y(n3534) );
  CLKINVX1 U2666 ( .A(n2417), .Y(n2756) );
  NOR2X1 U2667 ( .A(n1442), .B(n1378), .Y(n3532) );
  CLKINVX1 U2668 ( .A(n2754), .Y(n3533) );
  CLKNAND2X2 U2669 ( .A(n1378), .B(n1442), .Y(n2754) );
  MXI2X1 U2670 ( .A(n3535), .B(n3536), .S0(n366), .Y(n2999) );
  OAI21X1 U2671 ( .A0(n1290), .A1(n3537), .B0(n3538), .Y(n3536) );
  MXI2X1 U2672 ( .A(n3539), .B(n3540), .S0(n2623), .Y(n3538) );
  OAI21X1 U2673 ( .A0(n3537), .A1(n396), .B0(n3541), .Y(n3535) );
  MXI2X1 U2674 ( .A(n3540), .B(n3539), .S0(n2623), .Y(n3541) );
  CLKINVX1 U2675 ( .A(n2236), .Y(n2623) );
  NOR2X1 U2676 ( .A(n1481), .B(n1417), .Y(n3539) );
  CLKINVX1 U2677 ( .A(n2621), .Y(n3540) );
  CLKNAND2X2 U2678 ( .A(n1417), .B(n1481), .Y(n2621) );
  AOI21X1 U2679 ( .A0(n921), .A1(n1442), .B0(n864), .Y(n3525) );
  AOI21X1 U2680 ( .A0(n1139), .A1(n934), .B0(n957), .Y(n3524) );
  OAI222X1 U2681 ( .A0(n1441), .A1(n3542), .B0(n1143), .B1(n3543), .C0(n3544), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[200]) );
  XOR2X1 U2682 ( .A(n3177), .B(n3545), .Y(n3544) );
  XOR2X1 U2683 ( .A(n3005), .B(n3141), .Y(n3545) );
  MXI2X1 U2684 ( .A(n3546), .B(n3547), .S0(n373), .Y(n3141) );
  OAI21X1 U2685 ( .A0(n1250), .A1(n3548), .B0(n3549), .Y(n3547) );
  MXI2X1 U2686 ( .A(n3550), .B(n3551), .S0(n2764), .Y(n3549) );
  OAI21X1 U2687 ( .A0(n3548), .A1(n410), .B0(n3552), .Y(n3546) );
  MXI2X1 U2688 ( .A(n3551), .B(n3550), .S0(n2764), .Y(n3552) );
  CLKINVX1 U2689 ( .A(n3553), .Y(n2764) );
  NOR2X1 U2690 ( .A(n1441), .B(n1377), .Y(n3550) );
  CLKINVX1 U2691 ( .A(n2762), .Y(n3551) );
  CLKNAND2X2 U2692 ( .A(n1377), .B(n1441), .Y(n2762) );
  MXI2X1 U2693 ( .A(n3554), .B(n3555), .S0(n367), .Y(n3005) );
  OAI21X1 U2694 ( .A0(n1289), .A1(n3556), .B0(n3557), .Y(n3555) );
  MXI2X1 U2695 ( .A(n3558), .B(n3559), .S0(n2630), .Y(n3557) );
  OAI21X1 U2696 ( .A0(n3556), .A1(n397), .B0(n3560), .Y(n3554) );
  MXI2X1 U2697 ( .A(n3559), .B(n3558), .S0(n2630), .Y(n3560) );
  CLKINVX1 U2698 ( .A(n2242), .Y(n2630) );
  NOR2X1 U2699 ( .A(n1480), .B(n1416), .Y(n3558) );
  CLKINVX1 U2700 ( .A(n2628), .Y(n3559) );
  CLKNAND2X2 U2701 ( .A(n1416), .B(n1480), .Y(n2628) );
  AOI21X1 U2702 ( .A0(n921), .A1(n1441), .B0(n864), .Y(n3543) );
  AOI21X1 U2703 ( .A0(n1143), .A1(n934), .B0(n957), .Y(n3542) );
  OAI222X1 U2704 ( .A0(n877), .A1(n3561), .B0(n3562), .B1(n905), .C0(
        Inst_AEAD_u_input_n320), .C1(n856), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[1]) );
  XOR2X1 U2705 ( .A(n3563), .B(n2227), .Y(n3562) );
  MXI2X1 U2706 ( .A(n2684), .B(n3564), .S0(n1475), .Y(n2227) );
  XOR2X1 U2707 ( .A(n1347), .B(n380), .Y(n2684) );
  XOR2X1 U2708 ( .A(n2144), .B(n1924), .Y(n3563) );
  MXI2X1 U2709 ( .A(n2761), .B(n3553), .S0(n1441), .Y(n1924) );
  XOR2X1 U2710 ( .A(n1313), .B(n373), .Y(n2761) );
  MXI2X1 U2711 ( .A(n2883), .B(n3565), .S0(n1434), .Y(n2144) );
  CLKINVX1 U2712 ( .A(n2886), .Y(n3565) );
  XNOR2X1 U2713 ( .A(n1306), .B(n1498), .Y(n2883) );
  OAI222X1 U2714 ( .A0(n877), .A1(n3566), .B0(n902), .B1(n3567), .C0(n853), 
        .C1(n1718), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[19]) );
  XNOR2X1 U2715 ( .A(n2226), .B(n3568), .Y(n3567) );
  XOR2X1 U2716 ( .A(n2193), .B(n2128), .Y(n3568) );
  MXI2X1 U2717 ( .A(n2508), .B(n3309), .S0(n1493), .Y(n2128) );
  XOR2X1 U2718 ( .A(n1365), .B(n358), .Y(n2508) );
  MXI2X1 U2719 ( .A(n2786), .B(n3239), .S0(n1459), .Y(n2193) );
  XNOR2X1 U2720 ( .A(n1268), .B(n454), .Y(n3239) );
  XNOR2X1 U2721 ( .A(n1331), .B(n1523), .Y(n2786) );
  OAI222X1 U2722 ( .A0(n1440), .A1(n3569), .B0(n1147), .B1(n3570), .C0(n3571), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[199]) );
  XNOR2X1 U2723 ( .A(n3572), .B(n3573), .Y(n3571) );
  XNOR2X1 U2724 ( .A(n3153), .B(n3011), .Y(n3572) );
  MXI2X1 U2725 ( .A(n3574), .B(n3575), .S0(n369), .Y(n3011) );
  OAI21X1 U2726 ( .A0(n1288), .A1(n3576), .B0(n3577), .Y(n3575) );
  MXI2X1 U2727 ( .A(n3578), .B(n3579), .S0(n2637), .Y(n3577) );
  OAI21X1 U2728 ( .A0(n3576), .A1(n398), .B0(n3580), .Y(n3574) );
  MXI2X1 U2729 ( .A(n3579), .B(n3578), .S0(n2637), .Y(n3580) );
  CLKINVX1 U2730 ( .A(n2251), .Y(n2637) );
  NOR2X1 U2731 ( .A(n1479), .B(n1415), .Y(n3578) );
  CLKINVX1 U2732 ( .A(n2635), .Y(n3579) );
  CLKNAND2X2 U2733 ( .A(n1415), .B(n1479), .Y(n2635) );
  MXI2X1 U2734 ( .A(n3581), .B(n3582), .S0(n350), .Y(n3153) );
  OAI21X1 U2735 ( .A0(n1249), .A1(n3583), .B0(n3584), .Y(n3582) );
  MXI2X1 U2736 ( .A(n3585), .B(n3586), .S0(n2783), .Y(n3584) );
  OAI2B1X1 U2737 ( .A1N(n1249), .A0(n3583), .B0(n3587), .Y(n3581) );
  MXI2X1 U2738 ( .A(n3586), .B(n3585), .S0(n2783), .Y(n3587) );
  NOR2X1 U2739 ( .A(n1440), .B(n2785), .Y(n3585) );
  CLKINVX1 U2740 ( .A(n2780), .Y(n3586) );
  CLKNAND2X2 U2741 ( .A(n1440), .B(n2785), .Y(n2780) );
  AOI21X1 U2742 ( .A0(n921), .A1(n1440), .B0(n864), .Y(n3570) );
  AOI21X1 U2743 ( .A0(n1147), .A1(n934), .B0(n957), .Y(n3569) );
  OAI222X1 U2744 ( .A0(n1439), .A1(n3588), .B0(n1151), .B1(n3589), .C0(n3590), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[198]) );
  XNOR2X1 U2745 ( .A(n3591), .B(n3592), .Y(n3590) );
  XNOR2X1 U2746 ( .A(n3165), .B(n3017), .Y(n3591) );
  MXI2X1 U2747 ( .A(n3593), .B(n3594), .S0(n355), .Y(n3017) );
  OAI21X1 U2748 ( .A0(n1287), .A1(n3595), .B0(n3596), .Y(n3594) );
  MXI2X1 U2749 ( .A(n3597), .B(n3598), .S0(n2648), .Y(n3596) );
  OAI21X1 U2750 ( .A0(n3595), .A1(n399), .B0(n3599), .Y(n3593) );
  MXI2X1 U2751 ( .A(n3598), .B(n3597), .S0(n2648), .Y(n3599) );
  CLKINVX1 U2752 ( .A(n2256), .Y(n2648) );
  NOR2X1 U2753 ( .A(n1478), .B(n1414), .Y(n3597) );
  CLKINVX1 U2754 ( .A(n2646), .Y(n3598) );
  CLKNAND2X2 U2755 ( .A(n1414), .B(n1478), .Y(n2646) );
  MXI2X1 U2756 ( .A(n3600), .B(n3601), .S0(n1503), .Y(n3165) );
  OAI2B1X1 U2757 ( .A1N(n1248), .A0(n3602), .B0(n3603), .Y(n3601) );
  MXI2X1 U2758 ( .A(n3604), .B(n3605), .S0(n2423), .Y(n3603) );
  OAI21X1 U2759 ( .A0(n1248), .A1(n3602), .B0(n3606), .Y(n3600) );
  MXI2X1 U2760 ( .A(n3605), .B(n3604), .S0(n2423), .Y(n3606) );
  CLKINVX1 U2761 ( .A(n2798), .Y(n3604) );
  CLKNAND2X2 U2762 ( .A(n1439), .B(n2801), .Y(n2798) );
  NOR2X1 U2763 ( .A(n1439), .B(n2801), .Y(n3605) );
  AOI21X1 U2764 ( .A0(n921), .A1(n1439), .B0(n865), .Y(n3589) );
  AOI21X1 U2765 ( .A0(n1151), .A1(n934), .B0(n957), .Y(n3588) );
  OAI222X1 U2766 ( .A0(n1438), .A1(n3607), .B0(n1155), .B1(n3608), .C0(n3609), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[197]) );
  XNOR2X1 U2767 ( .A(n3610), .B(n3611), .Y(n3609) );
  XNOR2X1 U2768 ( .A(n3177), .B(n3027), .Y(n3610) );
  MXI2X1 U2769 ( .A(n3612), .B(n3613), .S0(n357), .Y(n3027) );
  OAI21X1 U2770 ( .A0(n1286), .A1(n3614), .B0(n3615), .Y(n3613) );
  MXI2X1 U2771 ( .A(n3616), .B(n3617), .S0(n2659), .Y(n3615) );
  OAI21X1 U2772 ( .A0(n3614), .A1(n400), .B0(n3618), .Y(n3612) );
  MXI2X1 U2773 ( .A(n3617), .B(n3616), .S0(n2659), .Y(n3618) );
  CLKINVX1 U2774 ( .A(n2261), .Y(n2659) );
  NOR2X1 U2775 ( .A(n1477), .B(n1413), .Y(n3616) );
  CLKINVX1 U2776 ( .A(n2657), .Y(n3617) );
  CLKNAND2X2 U2777 ( .A(n1413), .B(n1477), .Y(n2657) );
  MXI2X1 U2778 ( .A(n3619), .B(n3620), .S0(n1502), .Y(n3177) );
  OAI2B1X1 U2779 ( .A1N(n1247), .A0(n3621), .B0(n3622), .Y(n3620) );
  MXI2X1 U2780 ( .A(n3623), .B(n3624), .S0(n2491), .Y(n3622) );
  OAI21X1 U2781 ( .A0(n1247), .A1(n3621), .B0(n3625), .Y(n3619) );
  MXI2X1 U2782 ( .A(n3624), .B(n3623), .S0(n2491), .Y(n3625) );
  CLKINVX1 U2783 ( .A(n2814), .Y(n3623) );
  CLKNAND2X2 U2784 ( .A(n1438), .B(n2817), .Y(n2814) );
  NOR2X1 U2785 ( .A(n1438), .B(n2817), .Y(n3624) );
  AOI21X1 U2786 ( .A0(n921), .A1(n1438), .B0(n865), .Y(n3608) );
  AOI21X1 U2787 ( .A0(n1155), .A1(n934), .B0(n957), .Y(n3607) );
  OAI222X1 U2788 ( .A0(n1437), .A1(n3626), .B0(n1159), .B1(n3627), .C0(n3628), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[196]) );
  XNOR2X1 U2789 ( .A(n3629), .B(n3630), .Y(n3628) );
  XNOR2X1 U2790 ( .A(n3189), .B(n3033), .Y(n3629) );
  MX2X1 U2791 ( .A(n3631), .B(n3632), .S0(n1540), .Y(n3033) );
  OAI21X1 U2792 ( .A0(n3633), .A1(n401), .B0(n3634), .Y(n3632) );
  MXI2X1 U2793 ( .A(n3635), .B(n3636), .S0(n2674), .Y(n3634) );
  OAI21X1 U2794 ( .A0(n1285), .A1(n3633), .B0(n3637), .Y(n3631) );
  MXI2X1 U2795 ( .A(n3636), .B(n3635), .S0(n2674), .Y(n3637) );
  CLKINVX1 U2796 ( .A(n2415), .Y(n2674) );
  CLKINVX1 U2797 ( .A(n2672), .Y(n3635) );
  CLKNAND2X2 U2798 ( .A(n1412), .B(n1476), .Y(n2672) );
  NOR2X1 U2799 ( .A(n1476), .B(n1412), .Y(n3636) );
  CLKINVX1 U2800 ( .A(n3573), .Y(n3189) );
  MXI2X1 U2801 ( .A(n3638), .B(n3639), .S0(n1501), .Y(n3573) );
  OAI2B1X1 U2802 ( .A1N(n1246), .A0(n3640), .B0(n3641), .Y(n3639) );
  MXI2X1 U2803 ( .A(n3642), .B(n3643), .S0(n2590), .Y(n3641) );
  OAI21X1 U2804 ( .A0(n1246), .A1(n3640), .B0(n3644), .Y(n3638) );
  MXI2X1 U2805 ( .A(n3643), .B(n3642), .S0(n2590), .Y(n3644) );
  CLKINVX1 U2806 ( .A(n2830), .Y(n3642) );
  CLKNAND2X2 U2807 ( .A(n1437), .B(n2833), .Y(n2830) );
  NOR2X1 U2808 ( .A(n1437), .B(n2833), .Y(n3643) );
  AOI21X1 U2809 ( .A0(n921), .A1(n1437), .B0(n865), .Y(n3627) );
  AOI21X1 U2810 ( .A0(n1159), .A1(n934), .B0(n957), .Y(n3626) );
  OAI222X1 U2811 ( .A0(n1436), .A1(n3645), .B0(n1163), .B1(n3646), .C0(n3647), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[195]) );
  XNOR2X1 U2812 ( .A(n3648), .B(n3649), .Y(n3647) );
  XNOR2X1 U2813 ( .A(n3201), .B(n3039), .Y(n3648) );
  MX2X1 U2814 ( .A(n3650), .B(n3651), .S0(n1539), .Y(n3039) );
  OAI21X1 U2815 ( .A0(n3652), .A1(n402), .B0(n3653), .Y(n3651) );
  MXI2X1 U2816 ( .A(n3654), .B(n3655), .S0(n2687), .Y(n3653) );
  OAI21X1 U2817 ( .A0(n1284), .A1(n3652), .B0(n3656), .Y(n3650) );
  MXI2X1 U2818 ( .A(n3655), .B(n3654), .S0(n2687), .Y(n3656) );
  CLKINVX1 U2819 ( .A(n3564), .Y(n2687) );
  CLKINVX1 U2820 ( .A(n2685), .Y(n3654) );
  CLKNAND2X2 U2821 ( .A(n1411), .B(n1475), .Y(n2685) );
  NOR2X1 U2822 ( .A(n1475), .B(n1411), .Y(n3655) );
  CLKINVX1 U2823 ( .A(n3592), .Y(n3201) );
  MXI2X1 U2824 ( .A(n3657), .B(n3658), .S0(n1500), .Y(n3592) );
  OAI2B1X1 U2825 ( .A1N(n1245), .A0(n3659), .B0(n3660), .Y(n3658) );
  MXI2X1 U2826 ( .A(n3661), .B(n3662), .S0(n2699), .Y(n3660) );
  OAI21X1 U2827 ( .A0(n1245), .A1(n3659), .B0(n3663), .Y(n3657) );
  MXI2X1 U2828 ( .A(n3662), .B(n3661), .S0(n2699), .Y(n3663) );
  CLKINVX1 U2829 ( .A(n2853), .Y(n3661) );
  CLKNAND2X2 U2830 ( .A(n1436), .B(n2856), .Y(n2853) );
  NOR2X1 U2831 ( .A(n1436), .B(n2856), .Y(n3662) );
  AOI21X1 U2832 ( .A0(n921), .A1(n1436), .B0(n865), .Y(n3646) );
  AOI21X1 U2833 ( .A0(n1163), .A1(n934), .B0(n957), .Y(n3645) );
  OAI222X1 U2834 ( .A0(n1435), .A1(n3664), .B0(n1167), .B1(n3665), .C0(n3666), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[194]) );
  XNOR2X1 U2835 ( .A(n3218), .B(n3667), .Y(n3666) );
  XOR2X1 U2836 ( .A(n2921), .B(n3045), .Y(n3667) );
  MXI2X1 U2837 ( .A(n3668), .B(n3669), .S0(n370), .Y(n3045) );
  OAI21X1 U2838 ( .A0(n1283), .A1(n3670), .B0(n3671), .Y(n3669) );
  MXI2X1 U2839 ( .A(n3672), .B(n3673), .S0(n2707), .Y(n3671) );
  OAI21X1 U2840 ( .A0(n3670), .A1(n403), .B0(n3674), .Y(n3668) );
  MXI2X1 U2841 ( .A(n3673), .B(n3672), .S0(n2707), .Y(n3674) );
  CLKINVX1 U2842 ( .A(n3675), .Y(n2707) );
  NOR2X1 U2843 ( .A(n1474), .B(n1410), .Y(n3672) );
  CLKINVX1 U2844 ( .A(n2705), .Y(n3673) );
  CLKNAND2X2 U2845 ( .A(n1410), .B(n1474), .Y(n2705) );
  MXI2X1 U2846 ( .A(n3676), .B(n3677), .S0(n1560), .Y(n2921) );
  OAI21X1 U2847 ( .A0(n3678), .A1(n381), .B0(n3679), .Y(n3677) );
  MXI2X1 U2848 ( .A(n3680), .B(n3681), .S0(n2472), .Y(n3679) );
  OAI21X1 U2849 ( .A0(n1305), .A1(n3678), .B0(n3682), .Y(n3676) );
  MXI2X1 U2850 ( .A(n3681), .B(n3680), .S0(n2472), .Y(n3682) );
  CLKINVX1 U2851 ( .A(n3089), .Y(n2472) );
  CLKINVX1 U2852 ( .A(n2470), .Y(n3680) );
  CLKNAND2X2 U2853 ( .A(n1432), .B(n1496), .Y(n2470) );
  NOR2X1 U2854 ( .A(n1496), .B(n1432), .Y(n3681) );
  CLKINVX1 U2855 ( .A(n3611), .Y(n3218) );
  MXI2X1 U2856 ( .A(n3683), .B(n3684), .S0(n1499), .Y(n3611) );
  OAI2B1X1 U2857 ( .A1N(n1244), .A0(n3685), .B0(n3686), .Y(n3684) );
  MXI2X1 U2858 ( .A(n3687), .B(n3688), .S0(n2849), .Y(n3686) );
  OAI21X1 U2859 ( .A0(n1244), .A1(n3685), .B0(n3689), .Y(n3683) );
  MXI2X1 U2860 ( .A(n3688), .B(n3687), .S0(n2849), .Y(n3689) );
  CLKINVX1 U2861 ( .A(n2868), .Y(n3687) );
  CLKNAND2X2 U2862 ( .A(n1435), .B(n2871), .Y(n2868) );
  NOR2X1 U2863 ( .A(n1435), .B(n2871), .Y(n3688) );
  AOI21X1 U2864 ( .A0(n922), .A1(n1435), .B0(n865), .Y(n3665) );
  AOI21X1 U2865 ( .A0(n1167), .A1(n934), .B0(n957), .Y(n3664) );
  OAI222X1 U2866 ( .A0(n1434), .A1(n3690), .B0(n1171), .B1(n3691), .C0(n3692), 
        .C1(n896), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[193]) );
  XNOR2X1 U2867 ( .A(n3231), .B(n3693), .Y(n3692) );
  XOR2X1 U2868 ( .A(n2929), .B(n3051), .Y(n3693) );
  MXI2X1 U2869 ( .A(n3694), .B(n3695), .S0(n363), .Y(n3051) );
  OAI21X1 U2870 ( .A0(n1282), .A1(n3696), .B0(n3697), .Y(n3695) );
  MXI2X1 U2871 ( .A(n3698), .B(n3699), .S0(n2719), .Y(n3697) );
  OAI21X1 U2872 ( .A0(n3696), .A1(n404), .B0(n3700), .Y(n3694) );
  MXI2X1 U2873 ( .A(n3699), .B(n3698), .S0(n2719), .Y(n3700) );
  CLKINVX1 U2874 ( .A(n2275), .Y(n2719) );
  NOR2X1 U2875 ( .A(n1473), .B(n1409), .Y(n3698) );
  CLKINVX1 U2876 ( .A(n2717), .Y(n3699) );
  CLKNAND2X2 U2877 ( .A(n1409), .B(n1473), .Y(n2717) );
  MXI2X1 U2878 ( .A(n3701), .B(n3702), .S0(n354), .Y(n2929) );
  OAI21X1 U2879 ( .A0(n1304), .A1(n3703), .B0(n3704), .Y(n3702) );
  MXI2X1 U2880 ( .A(n3705), .B(n3706), .S0(n2482), .Y(n3704) );
  OAI21X1 U2881 ( .A0(n3703), .A1(n382), .B0(n3707), .Y(n3701) );
  MXI2X1 U2882 ( .A(n3706), .B(n3705), .S0(n2482), .Y(n3707) );
  CLKINVX1 U2883 ( .A(n3214), .Y(n2482) );
  NOR2X1 U2884 ( .A(n1495), .B(n1431), .Y(n3705) );
  CLKINVX1 U2885 ( .A(n2480), .Y(n3706) );
  CLKNAND2X2 U2886 ( .A(n1431), .B(n1495), .Y(n2480) );
  CLKINVX1 U2887 ( .A(n3630), .Y(n3231) );
  MXI2X1 U2888 ( .A(n3708), .B(n3709), .S0(n1498), .Y(n3630) );
  OAI2B1X1 U2889 ( .A1N(n1243), .A0(n3710), .B0(n3711), .Y(n3709) );
  MXI2X1 U2890 ( .A(n3712), .B(n3713), .S0(n2886), .Y(n3711) );
  OAI21X1 U2891 ( .A0(n1243), .A1(n3710), .B0(n3714), .Y(n3708) );
  MXI2X1 U2892 ( .A(n3713), .B(n3712), .S0(n2886), .Y(n3714) );
  CLKINVX1 U2893 ( .A(n2884), .Y(n3712) );
  CLKNAND2X2 U2894 ( .A(n1434), .B(n2888), .Y(n2884) );
  NOR2X1 U2895 ( .A(n1434), .B(n2888), .Y(n3713) );
  AOI21X1 U2896 ( .A0(n922), .A1(n1434), .B0(n865), .Y(n3691) );
  AOI21X1 U2897 ( .A0(n1171), .A1(n934), .B0(n957), .Y(n3690) );
  OAI222X1 U2898 ( .A0(n1433), .A1(n3715), .B0(n1175), .B1(n3716), .C0(n3717), 
        .C1(n897), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[192]) );
  XNOR2X1 U2899 ( .A(n3244), .B(n3718), .Y(n3717) );
  XOR2X1 U2900 ( .A(n2936), .B(n3057), .Y(n3718) );
  MXI2X1 U2901 ( .A(n3719), .B(n3720), .S0(n351), .Y(n3057) );
  OAI21X1 U2902 ( .A0(n1281), .A1(n3721), .B0(n3722), .Y(n3720) );
  MXI2X1 U2903 ( .A(n3723), .B(n2729), .S0(n2280), .Y(n3722) );
  OAI21X1 U2904 ( .A0(n3721), .A1(n411), .B0(n3724), .Y(n3719) );
  MXI2X1 U2905 ( .A(n2729), .B(n3723), .S0(n2280), .Y(n3724) );
  NOR2X1 U2906 ( .A(n1472), .B(n1408), .Y(n3723) );
  AND2X1 U2907 ( .A(n1408), .B(n1472), .Y(n2729) );
  MXI2X1 U2908 ( .A(n3725), .B(n3726), .S0(n356), .Y(n2936) );
  OAI21X1 U2909 ( .A0(n1303), .A1(n3727), .B0(n3728), .Y(n3726) );
  MXI2X1 U2910 ( .A(n3729), .B(n3730), .S0(n2501), .Y(n3728) );
  OAI21X1 U2911 ( .A0(n3727), .A1(n383), .B0(n3731), .Y(n3725) );
  MXI2X1 U2912 ( .A(n3730), .B(n3729), .S0(n2501), .Y(n3731) );
  CLKINVX1 U2913 ( .A(n3369), .Y(n2501) );
  NOR2X1 U2914 ( .A(n1494), .B(n1430), .Y(n3729) );
  CLKINVX1 U2915 ( .A(n2499), .Y(n3730) );
  CLKNAND2X2 U2916 ( .A(n1430), .B(n1494), .Y(n2499) );
  CLKINVX1 U2917 ( .A(n3649), .Y(n3244) );
  MXI2X1 U2918 ( .A(n3732), .B(n3733), .S0(n1497), .Y(n3649) );
  OAI21X1 U2919 ( .A0(n3734), .A1(n378), .B0(n3735), .Y(n3733) );
  MXI2X1 U2920 ( .A(n3736), .B(n3737), .S0(n2905), .Y(n3735) );
  OAI21X1 U2921 ( .A0(n1242), .A1(n3734), .B0(n3738), .Y(n3732) );
  MXI2X1 U2922 ( .A(n3737), .B(n3736), .S0(n2905), .Y(n3738) );
  CLKINVX1 U2923 ( .A(n2903), .Y(n3736) );
  CLKNAND2X2 U2924 ( .A(n1433), .B(n2907), .Y(n2903) );
  NOR2X1 U2925 ( .A(n1433), .B(n2907), .Y(n3737) );
  AOI21X1 U2926 ( .A0(n922), .A1(n1433), .B0(n865), .Y(n3716) );
  AOI21X1 U2927 ( .A0(n1175), .A1(n935), .B0(n956), .Y(n3715) );
  OAI222X1 U2928 ( .A0(n1432), .A1(n3739), .B0(n1050), .B1(n3740), .C0(n887), 
        .C1(n3741), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[191]) );
  XOR2X1 U2929 ( .A(n3742), .B(n3743), .Y(n3741) );
  XOR2X1 U2930 ( .A(n3744), .B(n3745), .Y(n3743) );
  AOI21X1 U2931 ( .A0(n922), .A1(n1432), .B0(n866), .Y(n3740) );
  AOI21X1 U2932 ( .A0(n1050), .A1(n935), .B0(n956), .Y(n3739) );
  OAI222X1 U2933 ( .A0(n1431), .A1(n3746), .B0(n1054), .B1(n3747), .C0(n888), 
        .C1(n3748), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[190]) );
  XOR2X1 U2934 ( .A(n3749), .B(n3750), .Y(n3748) );
  XNOR2X1 U2935 ( .A(n3751), .B(n3745), .Y(n3750) );
  AOI21X1 U2936 ( .A0(n922), .A1(n1431), .B0(n866), .Y(n3747) );
  AOI21X1 U2937 ( .A0(n1054), .A1(n935), .B0(n956), .Y(n3746) );
  OAI222X1 U2938 ( .A0(n877), .A1(n3752), .B0(n903), .B1(n3753), .C0(n853), 
        .C1(n1717), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[18]) );
  XOR2X1 U2939 ( .A(n2234), .B(n3754), .Y(n3753) );
  XOR2X1 U2940 ( .A(n2197), .B(n2139), .Y(n3754) );
  MXI2X1 U2941 ( .A(n2519), .B(n3327), .S0(n1492), .Y(n2139) );
  XOR2X1 U2942 ( .A(n1364), .B(n360), .Y(n2519) );
  MXI2X1 U2943 ( .A(n2802), .B(n3252), .S0(n1458), .Y(n2197) );
  XNOR2X1 U2944 ( .A(n1267), .B(n455), .Y(n3252) );
  XNOR2X1 U2945 ( .A(n1330), .B(n1522), .Y(n2802) );
  OAI222X1 U2946 ( .A0(n1430), .A1(n3755), .B0(n1058), .B1(n3756), .C0(n887), 
        .C1(n3757), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[189]) );
  XOR2X1 U2947 ( .A(n3758), .B(n3759), .Y(n3757) );
  XNOR2X1 U2948 ( .A(n3760), .B(n3751), .Y(n3759) );
  AOI21X1 U2949 ( .A0(n922), .A1(n1430), .B0(n866), .Y(n3756) );
  AOI21X1 U2950 ( .A0(n1058), .A1(n935), .B0(n956), .Y(n3755) );
  OAI222X1 U2951 ( .A0(n1429), .A1(n3761), .B0(n1062), .B1(n3762), .C0(n888), 
        .C1(n3763), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[188]) );
  XOR2X1 U2952 ( .A(n3764), .B(n3765), .Y(n3763) );
  XNOR2X1 U2953 ( .A(n3766), .B(n3760), .Y(n3765) );
  AOI21X1 U2954 ( .A0(n922), .A1(n1429), .B0(n866), .Y(n3762) );
  AOI21X1 U2955 ( .A0(n1062), .A1(n935), .B0(n956), .Y(n3761) );
  OAI222X1 U2956 ( .A0(n1428), .A1(n3767), .B0(n1066), .B1(n3768), .C0(n888), 
        .C1(n3769), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[187]) );
  XOR2X1 U2957 ( .A(n3770), .B(n3771), .Y(n3769) );
  XNOR2X1 U2958 ( .A(n3772), .B(n3766), .Y(n3771) );
  AOI21X1 U2959 ( .A0(n922), .A1(n1428), .B0(n866), .Y(n3768) );
  AOI21X1 U2960 ( .A0(n1066), .A1(n935), .B0(n956), .Y(n3767) );
  OAI222X1 U2961 ( .A0(n1427), .A1(n3773), .B0(n1070), .B1(n3774), .C0(n888), 
        .C1(n3775), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[186]) );
  XOR2X1 U2962 ( .A(n3776), .B(n3777), .Y(n3775) );
  XNOR2X1 U2963 ( .A(n3744), .B(n3772), .Y(n3777) );
  AOI21X1 U2964 ( .A0(n922), .A1(n1427), .B0(n866), .Y(n3774) );
  AOI21X1 U2965 ( .A0(n1070), .A1(n935), .B0(n956), .Y(n3773) );
  OAI222X1 U2966 ( .A0(n1426), .A1(n3778), .B0(n1074), .B1(n3779), .C0(n888), 
        .C1(n3780), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[185]) );
  XOR2X1 U2967 ( .A(n3781), .B(n3782), .Y(n3780) );
  XOR2X1 U2968 ( .A(n3745), .B(n3776), .Y(n3782) );
  XOR2X1 U2969 ( .A(n3783), .B(n3678), .Y(n3745) );
  CLKNAND2X2 U2970 ( .A(n1368), .B(n381), .Y(n3783) );
  AOI21X1 U2971 ( .A0(n922), .A1(n1426), .B0(n866), .Y(n3779) );
  AOI21X1 U2972 ( .A0(n1074), .A1(n935), .B0(n956), .Y(n3778) );
  OAI222X1 U2973 ( .A0(n1425), .A1(n3784), .B0(n1078), .B1(n3785), .C0(n888), 
        .C1(n3786), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[184]) );
  XOR2X1 U2974 ( .A(n3787), .B(n3788), .Y(n3786) );
  XOR2X1 U2975 ( .A(n3751), .B(n3781), .Y(n3788) );
  XOR2X1 U2976 ( .A(n3789), .B(n3703), .Y(n3751) );
  CLKINVX1 U2977 ( .A(n3790), .Y(n3703) );
  CLKNAND2X2 U2978 ( .A(n1367), .B(n382), .Y(n3789) );
  AOI21X1 U2979 ( .A0(n922), .A1(n1425), .B0(n866), .Y(n3785) );
  AOI21X1 U2980 ( .A0(n1078), .A1(n936), .B0(n956), .Y(n3784) );
  OAI222X1 U2981 ( .A0(n1424), .A1(n3791), .B0(n1082), .B1(n3792), .C0(n888), 
        .C1(n3793), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[183]) );
  XOR2X1 U2982 ( .A(n3794), .B(n3795), .Y(n3793) );
  XOR2X1 U2983 ( .A(n3760), .B(n3787), .Y(n3795) );
  XOR2X1 U2984 ( .A(n3796), .B(n3727), .Y(n3760) );
  CLKINVX1 U2985 ( .A(n3797), .Y(n3727) );
  CLKNAND2X2 U2986 ( .A(n1366), .B(n383), .Y(n3796) );
  AOI21X1 U2987 ( .A0(n922), .A1(n1424), .B0(n866), .Y(n3792) );
  AOI21X1 U2988 ( .A0(n1082), .A1(n936), .B0(n956), .Y(n3791) );
  OAI222X1 U2989 ( .A0(n1423), .A1(n3798), .B0(n1086), .B1(n3799), .C0(n888), 
        .C1(n3800), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[182]) );
  XOR2X1 U2990 ( .A(n3801), .B(n3802), .Y(n3800) );
  XOR2X1 U2991 ( .A(n3766), .B(n3794), .Y(n3802) );
  XOR2X1 U2992 ( .A(n3803), .B(n3304), .Y(n3766) );
  CLKINVX1 U2993 ( .A(n3804), .Y(n3304) );
  CLKNAND2X2 U2994 ( .A(n1365), .B(n384), .Y(n3803) );
  AOI21X1 U2995 ( .A0(n923), .A1(n1423), .B0(n866), .Y(n3799) );
  AOI21X1 U2996 ( .A0(n1086), .A1(n936), .B0(n956), .Y(n3798) );
  OAI222X1 U2997 ( .A0(n1422), .A1(n3805), .B0(n1090), .B1(n3806), .C0(n888), 
        .C1(n3807), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[181]) );
  XOR2X1 U2998 ( .A(n3808), .B(n3809), .Y(n3807) );
  XOR2X1 U2999 ( .A(n3772), .B(n3801), .Y(n3809) );
  XOR2X1 U3000 ( .A(n3810), .B(n3322), .Y(n3772) );
  CLKINVX1 U3001 ( .A(n3811), .Y(n3322) );
  CLKNAND2X2 U3002 ( .A(n1364), .B(n385), .Y(n3810) );
  AOI21X1 U3003 ( .A0(n923), .A1(n1422), .B0(n866), .Y(n3806) );
  AOI21X1 U3004 ( .A0(n1090), .A1(n936), .B0(n956), .Y(n3805) );
  OAI222X1 U3005 ( .A0(n1421), .A1(n3812), .B0(n1094), .B1(n3813), .C0(n888), 
        .C1(n3814), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[180]) );
  XOR2X1 U3006 ( .A(n3815), .B(n3816), .Y(n3814) );
  XOR2X1 U3007 ( .A(n3776), .B(n3808), .Y(n3816) );
  XOR2X1 U3008 ( .A(n3817), .B(n3340), .Y(n3776) );
  CLKNAND2X2 U3009 ( .A(n1363), .B(n386), .Y(n3817) );
  AOI21X1 U3010 ( .A0(n923), .A1(n1421), .B0(n866), .Y(n3813) );
  AOI21X1 U3011 ( .A0(n1094), .A1(n936), .B0(n956), .Y(n3812) );
  OAI222X1 U3012 ( .A0(n877), .A1(n3818), .B0(n902), .B1(n3819), .C0(n853), 
        .C1(n1716), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[17]) );
  XOR2X1 U3013 ( .A(n2239), .B(n3820), .Y(n3819) );
  XOR2X1 U3014 ( .A(n2201), .B(n2145), .Y(n3820) );
  MXI2X1 U3015 ( .A(n2528), .B(n3345), .S0(n1491), .Y(n2145) );
  XOR2X1 U3016 ( .A(n1363), .B(n362), .Y(n2528) );
  MXI2X1 U3017 ( .A(n2818), .B(n3264), .S0(n1457), .Y(n2201) );
  XNOR2X1 U3018 ( .A(n1266), .B(n456), .Y(n3264) );
  XNOR2X1 U3019 ( .A(n1329), .B(n1521), .Y(n2818) );
  OAI222X1 U3020 ( .A0(n1420), .A1(n3821), .B0(n1098), .B1(n3822), .C0(n888), 
        .C1(n3823), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[179]) );
  XOR2X1 U3021 ( .A(n3824), .B(n3825), .Y(n3823) );
  XOR2X1 U3022 ( .A(n3781), .B(n3815), .Y(n3825) );
  XOR2X1 U3023 ( .A(n3826), .B(n3360), .Y(n3781) );
  CLKNAND2X2 U3024 ( .A(n1362), .B(n387), .Y(n3826) );
  AOI21X1 U3025 ( .A0(n923), .A1(n1420), .B0(n866), .Y(n3822) );
  AOI21X1 U3026 ( .A0(n1098), .A1(n936), .B0(n955), .Y(n3821) );
  OAI222X1 U3027 ( .A0(n1419), .A1(n3827), .B0(n1102), .B1(n3828), .C0(n888), 
        .C1(n3829), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[178]) );
  XOR2X1 U3028 ( .A(n3830), .B(n3831), .Y(n3829) );
  XOR2X1 U3029 ( .A(n3787), .B(n3824), .Y(n3831) );
  XOR2X1 U3030 ( .A(n3832), .B(n3384), .Y(n3787) );
  CLKNAND2X2 U3031 ( .A(n1361), .B(n388), .Y(n3832) );
  AOI21X1 U3032 ( .A0(n923), .A1(n1419), .B0(n866), .Y(n3828) );
  AOI21X1 U3033 ( .A0(n1102), .A1(n936), .B0(n955), .Y(n3827) );
  OAI222X1 U3034 ( .A0(n1418), .A1(n3833), .B0(n1106), .B1(n3834), .C0(n888), 
        .C1(n3835), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[177]) );
  XOR2X1 U3035 ( .A(n3836), .B(n3837), .Y(n3835) );
  XOR2X1 U3036 ( .A(n3794), .B(n3830), .Y(n3837) );
  XOR2X1 U3037 ( .A(n3838), .B(n3404), .Y(n3794) );
  CLKNAND2X2 U3038 ( .A(n1360), .B(n389), .Y(n3838) );
  AOI21X1 U3039 ( .A0(n923), .A1(n1418), .B0(n866), .Y(n3834) );
  AOI21X1 U3040 ( .A0(n1106), .A1(n936), .B0(n955), .Y(n3833) );
  OAI222X1 U3041 ( .A0(n1417), .A1(n3839), .B0(n1110), .B1(n3840), .C0(n889), 
        .C1(n3841), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[176]) );
  XOR2X1 U3042 ( .A(n3842), .B(n3843), .Y(n3841) );
  XOR2X1 U3043 ( .A(n3801), .B(n3836), .Y(n3843) );
  XOR2X1 U3044 ( .A(n3844), .B(n3424), .Y(n3801) );
  CLKNAND2X2 U3045 ( .A(n1359), .B(n390), .Y(n3844) );
  AOI21X1 U3046 ( .A0(n923), .A1(n1417), .B0(n866), .Y(n3840) );
  AOI21X1 U3047 ( .A0(n1110), .A1(n936), .B0(n955), .Y(n3839) );
  OAI222X1 U3048 ( .A0(n1416), .A1(n3845), .B0(n1114), .B1(n3846), .C0(n889), 
        .C1(n3847), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[175]) );
  XOR2X1 U3049 ( .A(n3848), .B(n3849), .Y(n3847) );
  XOR2X1 U3050 ( .A(n3808), .B(n3842), .Y(n3849) );
  XOR2X1 U3051 ( .A(n3850), .B(n3444), .Y(n3808) );
  CLKNAND2X2 U3052 ( .A(n1358), .B(n391), .Y(n3850) );
  AOI21X1 U3053 ( .A0(n923), .A1(n1416), .B0(n866), .Y(n3846) );
  AOI21X1 U3054 ( .A0(n1114), .A1(n920), .B0(n955), .Y(n3845) );
  OAI222X1 U3055 ( .A0(n1415), .A1(n3851), .B0(n1118), .B1(n3852), .C0(n889), 
        .C1(n3853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[174]) );
  XOR2X1 U3056 ( .A(n3854), .B(n3855), .Y(n3853) );
  XOR2X1 U3057 ( .A(n3815), .B(n3848), .Y(n3855) );
  XNOR2X1 U3058 ( .A(n3856), .B(n3857), .Y(n3815) );
  CLKNAND2X2 U3059 ( .A(n1357), .B(n392), .Y(n3856) );
  AOI21X1 U3060 ( .A0(n923), .A1(n1415), .B0(n866), .Y(n3852) );
  AOI21X1 U3061 ( .A0(n1118), .A1(n923), .B0(n955), .Y(n3851) );
  OAI222X1 U3062 ( .A0(n1414), .A1(n3858), .B0(n1122), .B1(n3859), .C0(n889), 
        .C1(n3860), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[173]) );
  XOR2X1 U3063 ( .A(n3861), .B(n3862), .Y(n3860) );
  XOR2X1 U3064 ( .A(n3824), .B(n3854), .Y(n3862) );
  XNOR2X1 U3065 ( .A(n3863), .B(n3864), .Y(n3824) );
  CLKNAND2X2 U3066 ( .A(n1356), .B(n393), .Y(n3863) );
  AOI21X1 U3067 ( .A0(n923), .A1(n1414), .B0(n866), .Y(n3859) );
  AOI21X1 U3068 ( .A0(n1122), .A1(n921), .B0(n955), .Y(n3858) );
  OAI222X1 U3069 ( .A0(n1413), .A1(n3865), .B0(n1126), .B1(n3866), .C0(n889), 
        .C1(n3867), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[172]) );
  XOR2X1 U3070 ( .A(n3868), .B(n3869), .Y(n3867) );
  XOR2X1 U3071 ( .A(n3830), .B(n3861), .Y(n3869) );
  XNOR2X1 U3072 ( .A(n3870), .B(n3871), .Y(n3830) );
  CLKNAND2X2 U3073 ( .A(n1355), .B(n394), .Y(n3870) );
  AOI21X1 U3074 ( .A0(n923), .A1(n1413), .B0(n866), .Y(n3866) );
  AOI21X1 U3075 ( .A0(n1126), .A1(n925), .B0(n955), .Y(n3865) );
  OAI222X1 U3076 ( .A0(n1412), .A1(n3872), .B0(n1130), .B1(n3873), .C0(n889), 
        .C1(n3874), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[171]) );
  XOR2X1 U3077 ( .A(n3875), .B(n3876), .Y(n3874) );
  XOR2X1 U3078 ( .A(n3836), .B(n3868), .Y(n3876) );
  XNOR2X1 U3079 ( .A(n3877), .B(n3878), .Y(n3836) );
  CLKNAND2X2 U3080 ( .A(n1354), .B(n395), .Y(n3877) );
  AOI21X1 U3081 ( .A0(n923), .A1(n1412), .B0(n866), .Y(n3873) );
  AOI21X1 U3082 ( .A0(n1130), .A1(n926), .B0(n955), .Y(n3872) );
  OAI222X1 U3083 ( .A0(n1411), .A1(n3879), .B0(n1134), .B1(n3880), .C0(n889), 
        .C1(n3881), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[170]) );
  XOR2X1 U3084 ( .A(n3882), .B(n3883), .Y(n3881) );
  XOR2X1 U3085 ( .A(n3842), .B(n3875), .Y(n3883) );
  XNOR2X1 U3086 ( .A(n3884), .B(n3885), .Y(n3842) );
  CLKNAND2X2 U3087 ( .A(n1353), .B(n396), .Y(n3884) );
  AOI21X1 U3088 ( .A0(n924), .A1(n1411), .B0(n866), .Y(n3880) );
  AOI21X1 U3089 ( .A0(n1134), .A1(n928), .B0(n955), .Y(n3879) );
  OAI222X1 U3090 ( .A0(n877), .A1(n3886), .B0(n902), .B1(n3887), .C0(n854), 
        .C1(n1715), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[16]) );
  XOR2X1 U3091 ( .A(n2205), .B(n3888), .Y(n3887) );
  XOR2X1 U3092 ( .A(n1860), .B(n2150), .Y(n3888) );
  MXI2X1 U3093 ( .A(n2537), .B(n3365), .S0(n1490), .Y(n2150) );
  XOR2X1 U3094 ( .A(n1362), .B(n344), .Y(n2537) );
  MXI2X1 U3095 ( .A(n2661), .B(n3401), .S0(n1449), .Y(n1860) );
  XOR2X1 U3096 ( .A(n1321), .B(n348), .Y(n2661) );
  MXI2X1 U3097 ( .A(n2834), .B(n3276), .S0(n1456), .Y(n2205) );
  XNOR2X1 U3098 ( .A(n1265), .B(n457), .Y(n3276) );
  XNOR2X1 U3099 ( .A(n1328), .B(n1520), .Y(n2834) );
  OAI222X1 U3100 ( .A0(n1410), .A1(n3889), .B0(n1138), .B1(n3890), .C0(n889), 
        .C1(n3891), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[169]) );
  XOR2X1 U3101 ( .A(n3892), .B(n3893), .Y(n3891) );
  XOR2X1 U3102 ( .A(n3848), .B(n3882), .Y(n3893) );
  XNOR2X1 U3103 ( .A(n3894), .B(n3895), .Y(n3848) );
  CLKNAND2X2 U3104 ( .A(n1352), .B(n397), .Y(n3894) );
  AOI21X1 U3105 ( .A0(n924), .A1(n1410), .B0(n866), .Y(n3890) );
  AOI21X1 U3106 ( .A0(n1138), .A1(n922), .B0(n955), .Y(n3889) );
  OAI222X1 U3107 ( .A0(n1409), .A1(n3896), .B0(n1142), .B1(n3897), .C0(n889), 
        .C1(n3898), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[168]) );
  XOR2X1 U3108 ( .A(n3899), .B(n3900), .Y(n3898) );
  XOR2X1 U3109 ( .A(n3854), .B(n3892), .Y(n3900) );
  XNOR2X1 U3110 ( .A(n3901), .B(n3902), .Y(n3854) );
  CLKNAND2X2 U3111 ( .A(n1351), .B(n398), .Y(n3901) );
  AOI21X1 U3112 ( .A0(n924), .A1(n1409), .B0(n866), .Y(n3897) );
  AOI21X1 U3113 ( .A0(n1142), .A1(n924), .B0(n955), .Y(n3896) );
  OAI222X1 U3114 ( .A0(n1408), .A1(n3903), .B0(n1146), .B1(n3904), .C0(n889), 
        .C1(n3905), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[167]) );
  XOR2X1 U3115 ( .A(n3906), .B(n3907), .Y(n3905) );
  XOR2X1 U3116 ( .A(n3861), .B(n3899), .Y(n3907) );
  XNOR2X1 U3117 ( .A(n3908), .B(n3909), .Y(n3861) );
  CLKNAND2X2 U3118 ( .A(n1350), .B(n399), .Y(n3908) );
  AOI21X1 U3119 ( .A0(n924), .A1(n1408), .B0(n866), .Y(n3904) );
  AOI21X1 U3120 ( .A0(n1146), .A1(n936), .B0(n955), .Y(n3903) );
  OAI222X1 U3121 ( .A0(n1407), .A1(n3910), .B0(n1150), .B1(n3911), .C0(n889), 
        .C1(n3912), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[166]) );
  XOR2X1 U3122 ( .A(n3913), .B(n3914), .Y(n3912) );
  XOR2X1 U3123 ( .A(n3868), .B(n3906), .Y(n3914) );
  XNOR2X1 U3124 ( .A(n3915), .B(n3916), .Y(n3868) );
  CLKNAND2X2 U3125 ( .A(n1349), .B(n400), .Y(n3915) );
  AOI21X1 U3126 ( .A0(n924), .A1(n1407), .B0(n867), .Y(n3911) );
  AOI21X1 U3127 ( .A0(n1150), .A1(n936), .B0(n954), .Y(n3910) );
  OAI222X1 U3128 ( .A0(n1406), .A1(n3917), .B0(n1154), .B1(n3918), .C0(n889), 
        .C1(n3919), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[165]) );
  XOR2X1 U3129 ( .A(n3920), .B(n3921), .Y(n3919) );
  XOR2X1 U3130 ( .A(n3875), .B(n3913), .Y(n3921) );
  XNOR2X1 U3131 ( .A(n3922), .B(n3923), .Y(n3875) );
  CLKNAND2X2 U3132 ( .A(n1348), .B(n401), .Y(n3922) );
  AOI21X1 U3133 ( .A0(n925), .A1(n1406), .B0(n867), .Y(n3918) );
  AOI21X1 U3134 ( .A0(n1154), .A1(n936), .B0(n954), .Y(n3917) );
  OAI222X1 U3135 ( .A0(n1405), .A1(n3924), .B0(n1158), .B1(n3925), .C0(n890), 
        .C1(n3926), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[164]) );
  XOR2X1 U3136 ( .A(n3927), .B(n3928), .Y(n3926) );
  XOR2X1 U3137 ( .A(n3882), .B(n3920), .Y(n3928) );
  XNOR2X1 U3138 ( .A(n3929), .B(n3930), .Y(n3882) );
  CLKNAND2X2 U3139 ( .A(n1347), .B(n402), .Y(n3929) );
  AOI21X1 U3140 ( .A0(n925), .A1(n1405), .B0(n867), .Y(n3925) );
  AOI21X1 U3141 ( .A0(n1158), .A1(n936), .B0(n954), .Y(n3924) );
  OAI222X1 U3142 ( .A0(n1404), .A1(n3931), .B0(n1162), .B1(n3932), .C0(n890), 
        .C1(n3933), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[163]) );
  XOR2X1 U3143 ( .A(n3934), .B(n3935), .Y(n3933) );
  XOR2X1 U3144 ( .A(n3892), .B(n3927), .Y(n3935) );
  XNOR2X1 U3145 ( .A(n3936), .B(n3937), .Y(n3892) );
  CLKNAND2X2 U3146 ( .A(n1346), .B(n403), .Y(n3936) );
  AOI21X1 U3147 ( .A0(n925), .A1(n1404), .B0(n867), .Y(n3932) );
  AOI21X1 U3148 ( .A0(n1162), .A1(n935), .B0(n954), .Y(n3931) );
  OAI222X1 U3149 ( .A0(n1403), .A1(n3938), .B0(n1166), .B1(n3939), .C0(n890), 
        .C1(n3940), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[162]) );
  XOR2X1 U3150 ( .A(n3941), .B(n3942), .Y(n3940) );
  XOR2X1 U3151 ( .A(n3899), .B(n3934), .Y(n3942) );
  XNOR2X1 U3152 ( .A(n3943), .B(n3944), .Y(n3899) );
  CLKNAND2X2 U3153 ( .A(n1345), .B(n404), .Y(n3943) );
  AOI21X1 U3154 ( .A0(n925), .A1(n1403), .B0(n867), .Y(n3939) );
  AOI21X1 U3155 ( .A0(n1166), .A1(n935), .B0(n954), .Y(n3938) );
  OAI222X1 U3156 ( .A0(n1402), .A1(n3945), .B0(n1170), .B1(n3946), .C0(n890), 
        .C1(n3947), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[161]) );
  XOR2X1 U3157 ( .A(n3948), .B(n3949), .Y(n3947) );
  XOR2X1 U3158 ( .A(n3906), .B(n3941), .Y(n3949) );
  XNOR2X1 U3159 ( .A(n3950), .B(n3951), .Y(n3906) );
  CLKNAND2X2 U3160 ( .A(n1344), .B(n411), .Y(n3950) );
  AOI21X1 U3161 ( .A0(n925), .A1(n1402), .B0(n867), .Y(n3946) );
  AOI21X1 U3162 ( .A0(n1170), .A1(n935), .B0(n954), .Y(n3945) );
  OAI222X1 U3163 ( .A0(n1401), .A1(n3952), .B0(n1174), .B1(n3953), .C0(n890), 
        .C1(n3954), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[160]) );
  XOR2X1 U3164 ( .A(n3955), .B(n3956), .Y(n3954) );
  XOR2X1 U3165 ( .A(n3913), .B(n3948), .Y(n3956) );
  XNOR2X1 U3166 ( .A(n3957), .B(n3958), .Y(n3913) );
  CLKNAND2X2 U3167 ( .A(n1343), .B(n412), .Y(n3957) );
  AOI21X1 U3168 ( .A0(n926), .A1(n1401), .B0(n867), .Y(n3953) );
  AOI21X1 U3169 ( .A0(n1174), .A1(n935), .B0(n954), .Y(n3952) );
  OAI222X1 U3170 ( .A0(n878), .A1(n3959), .B0(n902), .B1(n3960), .C0(n853), 
        .C1(n2669), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[15]) );
  XOR2X1 U3171 ( .A(n2210), .B(n3961), .Y(n3960) );
  XOR2X1 U3172 ( .A(n1923), .B(n2154), .Y(n3961) );
  MXI2X1 U3173 ( .A(n2546), .B(n3389), .S0(n1489), .Y(n2154) );
  XOR2X1 U3174 ( .A(n1361), .B(n345), .Y(n2546) );
  MXI2X1 U3175 ( .A(n2676), .B(n3421), .S0(n1448), .Y(n1923) );
  XOR2X1 U3176 ( .A(n1320), .B(n349), .Y(n2676) );
  MXI2X1 U3177 ( .A(n2857), .B(n3288), .S0(n1455), .Y(n2210) );
  XNOR2X1 U3178 ( .A(n1264), .B(n458), .Y(n3288) );
  XNOR2X1 U3179 ( .A(n1327), .B(n1519), .Y(n2857) );
  OAI222X1 U3180 ( .A0(n1400), .A1(n3962), .B0(n1049), .B1(n3963), .C0(n890), 
        .C1(n3964), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[159]) );
  XOR2X1 U3181 ( .A(n3965), .B(n3966), .Y(n3964) );
  XOR2X1 U3182 ( .A(n3920), .B(n3955), .Y(n3966) );
  XNOR2X1 U3183 ( .A(n3967), .B(n3968), .Y(n3920) );
  CLKNAND2X2 U3184 ( .A(n1342), .B(n413), .Y(n3967) );
  AOI21X1 U3185 ( .A0(n925), .A1(n1400), .B0(n867), .Y(n3963) );
  AOI21X1 U3186 ( .A0(n1049), .A1(n935), .B0(n954), .Y(n3962) );
  OAI222X1 U3187 ( .A0(n1399), .A1(n3969), .B0(n1053), .B1(n3970), .C0(n890), 
        .C1(n3971), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[158]) );
  XOR2X1 U3188 ( .A(n3972), .B(n3973), .Y(n3971) );
  XOR2X1 U3189 ( .A(n3927), .B(n3965), .Y(n3973) );
  XNOR2X1 U3190 ( .A(n3974), .B(n3975), .Y(n3927) );
  CLKNAND2X2 U3191 ( .A(n1341), .B(n405), .Y(n3974) );
  AOI21X1 U3192 ( .A0(n926), .A1(n1399), .B0(n867), .Y(n3970) );
  AOI21X1 U3193 ( .A0(n1053), .A1(n934), .B0(n954), .Y(n3969) );
  OAI222X1 U3194 ( .A0(n1398), .A1(n3976), .B0(n1057), .B1(n3977), .C0(n890), 
        .C1(n3978), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[157]) );
  XOR2X1 U3195 ( .A(n3979), .B(n3980), .Y(n3978) );
  XOR2X1 U3196 ( .A(n3934), .B(n3972), .Y(n3980) );
  XNOR2X1 U3197 ( .A(n3981), .B(n3125), .Y(n3934) );
  XOR2X1 U3198 ( .A(n1404), .B(n1468), .Y(n3125) );
  CLKNAND2X2 U3199 ( .A(n1340), .B(n414), .Y(n3981) );
  AOI21X1 U3200 ( .A0(n926), .A1(n1398), .B0(n867), .Y(n3977) );
  AOI21X1 U3201 ( .A0(n1057), .A1(n934), .B0(n954), .Y(n3976) );
  OAI222X1 U3202 ( .A0(n1397), .A1(n3982), .B0(n1061), .B1(n3983), .C0(n890), 
        .C1(n3984), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[156]) );
  XOR2X1 U3203 ( .A(n3985), .B(n3986), .Y(n3984) );
  XOR2X1 U3204 ( .A(n3941), .B(n3979), .Y(n3986) );
  XNOR2X1 U3205 ( .A(n3987), .B(n3137), .Y(n3941) );
  XOR2X1 U3206 ( .A(n1403), .B(n1467), .Y(n3137) );
  CLKNAND2X2 U3207 ( .A(n1339), .B(n415), .Y(n3987) );
  AOI21X1 U3208 ( .A0(n926), .A1(n1397), .B0(n867), .Y(n3983) );
  AOI21X1 U3209 ( .A0(n1061), .A1(n934), .B0(n954), .Y(n3982) );
  OAI222X1 U3210 ( .A0(n1396), .A1(n3988), .B0(n1065), .B1(n3989), .C0(n890), 
        .C1(n3990), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[155]) );
  XOR2X1 U3211 ( .A(n3991), .B(n3992), .Y(n3990) );
  XOR2X1 U3212 ( .A(n3948), .B(n3985), .Y(n3992) );
  XNOR2X1 U3213 ( .A(n3993), .B(n3149), .Y(n3948) );
  XOR2X1 U3214 ( .A(n1402), .B(n1466), .Y(n3149) );
  CLKNAND2X2 U3215 ( .A(n1338), .B(n416), .Y(n3993) );
  AOI21X1 U3216 ( .A0(n926), .A1(n1396), .B0(n867), .Y(n3989) );
  AOI21X1 U3217 ( .A0(n1065), .A1(n934), .B0(n954), .Y(n3988) );
  OAI222X1 U3218 ( .A0(n1395), .A1(n3994), .B0(n1069), .B1(n3995), .C0(n890), 
        .C1(n3996), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[154]) );
  XOR2X1 U3219 ( .A(n3997), .B(n3998), .Y(n3996) );
  XOR2X1 U3220 ( .A(n3955), .B(n3991), .Y(n3998) );
  XNOR2X1 U3221 ( .A(n3999), .B(n3161), .Y(n3955) );
  XOR2X1 U3222 ( .A(n1401), .B(n1465), .Y(n3161) );
  CLKNAND2X2 U3223 ( .A(n1337), .B(n417), .Y(n3999) );
  AOI21X1 U3224 ( .A0(n926), .A1(n1395), .B0(n867), .Y(n3995) );
  AOI21X1 U3225 ( .A0(n1069), .A1(n933), .B0(n954), .Y(n3994) );
  OAI222X1 U3226 ( .A0(n1394), .A1(n4000), .B0(n1073), .B1(n4001), .C0(n890), 
        .C1(n4002), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[153]) );
  XOR2X1 U3227 ( .A(n4003), .B(n4004), .Y(n4002) );
  XOR2X1 U3228 ( .A(n3965), .B(n3997), .Y(n4004) );
  XNOR2X1 U3229 ( .A(n4005), .B(n3173), .Y(n3965) );
  XOR2X1 U3230 ( .A(n1400), .B(n1464), .Y(n3173) );
  CLKNAND2X2 U3231 ( .A(n1336), .B(n418), .Y(n4005) );
  AOI21X1 U3232 ( .A0(n926), .A1(n1394), .B0(n867), .Y(n4001) );
  AOI21X1 U3233 ( .A0(n1073), .A1(n933), .B0(n953), .Y(n4000) );
  OAI222X1 U3234 ( .A0(n1393), .A1(n4006), .B0(n1077), .B1(n4007), .C0(n890), 
        .C1(n4008), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[152]) );
  XOR2X1 U3235 ( .A(n4009), .B(n4010), .Y(n4008) );
  XOR2X1 U3236 ( .A(n3972), .B(n4003), .Y(n4010) );
  XNOR2X1 U3237 ( .A(n4011), .B(n3185), .Y(n3972) );
  XOR2X1 U3238 ( .A(n1399), .B(n1463), .Y(n3185) );
  CLKNAND2X2 U3239 ( .A(n1335), .B(n419), .Y(n4011) );
  AOI21X1 U3240 ( .A0(n926), .A1(n1393), .B0(n867), .Y(n4007) );
  AOI21X1 U3241 ( .A0(n1077), .A1(n933), .B0(n953), .Y(n4006) );
  OAI222X1 U3242 ( .A0(n1392), .A1(n4012), .B0(n1081), .B1(n4013), .C0(n891), 
        .C1(n4014), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[151]) );
  XOR2X1 U3243 ( .A(n4015), .B(n4016), .Y(n4014) );
  XOR2X1 U3244 ( .A(n3979), .B(n4009), .Y(n4016) );
  XNOR2X1 U3245 ( .A(n4017), .B(n3197), .Y(n3979) );
  XOR2X1 U3246 ( .A(n1398), .B(n1462), .Y(n3197) );
  CLKNAND2X2 U3247 ( .A(n1334), .B(n420), .Y(n4017) );
  AOI21X1 U3248 ( .A0(n927), .A1(n1392), .B0(n867), .Y(n4013) );
  AOI21X1 U3249 ( .A0(n1081), .A1(n933), .B0(n953), .Y(n4012) );
  OAI222X1 U3250 ( .A0(n1391), .A1(n4018), .B0(n1085), .B1(n4019), .C0(n891), 
        .C1(n4020), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[150]) );
  XOR2X1 U3251 ( .A(n4021), .B(n4022), .Y(n4020) );
  XOR2X1 U3252 ( .A(n3985), .B(n4015), .Y(n4022) );
  XNOR2X1 U3253 ( .A(n4023), .B(n3210), .Y(n3985) );
  XOR2X1 U3254 ( .A(n1397), .B(n1461), .Y(n3210) );
  CLKNAND2X2 U3255 ( .A(n1333), .B(n421), .Y(n4023) );
  AOI21X1 U3256 ( .A0(n925), .A1(n1391), .B0(n867), .Y(n4019) );
  AOI21X1 U3257 ( .A0(n1085), .A1(n932), .B0(n953), .Y(n4018) );
  OAI222X1 U3258 ( .A0(n878), .A1(n4024), .B0(n903), .B1(n4025), .C0(
        Inst_AEAD_u_input_n308), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[14]) );
  XOR2X1 U3259 ( .A(n2213), .B(n4026), .Y(n4025) );
  XOR2X1 U3260 ( .A(n2159), .B(n1980), .Y(n4026) );
  MXI2X1 U3261 ( .A(n2689), .B(n3441), .S0(n1447), .Y(n1980) );
  XOR2X1 U3262 ( .A(n1319), .B(n371), .Y(n2689) );
  MXI2X1 U3263 ( .A(n2554), .B(n3409), .S0(n1488), .Y(n2159) );
  XOR2X1 U3264 ( .A(n1360), .B(n346), .Y(n2554) );
  MXI2X1 U3265 ( .A(n2872), .B(n3300), .S0(n1454), .Y(n2213) );
  XNOR2X1 U3266 ( .A(n1263), .B(n459), .Y(n3300) );
  XNOR2X1 U3267 ( .A(n1326), .B(n1518), .Y(n2872) );
  OAI222X1 U3268 ( .A0(n1390), .A1(n4027), .B0(n1089), .B1(n4028), .C0(n891), 
        .C1(n4029), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[149]) );
  XOR2X1 U3269 ( .A(n4030), .B(n4031), .Y(n4029) );
  XOR2X1 U3270 ( .A(n3991), .B(n4021), .Y(n4031) );
  XNOR2X1 U3271 ( .A(n4032), .B(n3227), .Y(n3991) );
  XOR2X1 U3272 ( .A(n1396), .B(n1460), .Y(n3227) );
  CLKNAND2X2 U3273 ( .A(n1332), .B(n422), .Y(n4032) );
  AOI21X1 U3274 ( .A0(n927), .A1(n1390), .B0(n867), .Y(n4028) );
  AOI21X1 U3275 ( .A0(n1089), .A1(n932), .B0(n953), .Y(n4027) );
  OAI222X1 U3276 ( .A0(n1389), .A1(n4033), .B0(n1093), .B1(n4034), .C0(n891), 
        .C1(n4035), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[148]) );
  XOR2X1 U3277 ( .A(n4036), .B(n4037), .Y(n4035) );
  XOR2X1 U3278 ( .A(n3997), .B(n4030), .Y(n4037) );
  XNOR2X1 U3279 ( .A(n4038), .B(n3240), .Y(n3997) );
  XOR2X1 U3280 ( .A(n1395), .B(n1459), .Y(n3240) );
  CLKNAND2X2 U3281 ( .A(n1331), .B(n423), .Y(n4038) );
  AOI21X1 U3282 ( .A0(n927), .A1(n1389), .B0(n867), .Y(n4034) );
  AOI21X1 U3283 ( .A0(n1093), .A1(n932), .B0(n953), .Y(n4033) );
  OAI222X1 U3284 ( .A0(n1388), .A1(n4039), .B0(n1097), .B1(n4040), .C0(n891), 
        .C1(n4041), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[147]) );
  XOR2X1 U3285 ( .A(n4042), .B(n4043), .Y(n4041) );
  XOR2X1 U3286 ( .A(n4003), .B(n4036), .Y(n4043) );
  XNOR2X1 U3287 ( .A(n4044), .B(n3253), .Y(n4003) );
  XOR2X1 U3288 ( .A(n1394), .B(n1458), .Y(n3253) );
  CLKNAND2X2 U3289 ( .A(n1330), .B(n424), .Y(n4044) );
  AOI21X1 U3290 ( .A0(n927), .A1(n1388), .B0(n867), .Y(n4040) );
  AOI21X1 U3291 ( .A0(n1097), .A1(n932), .B0(n953), .Y(n4039) );
  OAI222X1 U3292 ( .A0(n1387), .A1(n4045), .B0(n1101), .B1(n4046), .C0(n891), 
        .C1(n4047), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[146]) );
  XOR2X1 U3293 ( .A(n4048), .B(n4049), .Y(n4047) );
  XOR2X1 U3294 ( .A(n4009), .B(n4042), .Y(n4049) );
  XNOR2X1 U3295 ( .A(n4050), .B(n3265), .Y(n4009) );
  XOR2X1 U3296 ( .A(n1393), .B(n1457), .Y(n3265) );
  CLKNAND2X2 U3297 ( .A(n1329), .B(n425), .Y(n4050) );
  AOI21X1 U3298 ( .A0(n927), .A1(n1387), .B0(n867), .Y(n4046) );
  AOI21X1 U3299 ( .A0(n1101), .A1(n932), .B0(n953), .Y(n4045) );
  OAI222X1 U3300 ( .A0(n1386), .A1(n4051), .B0(n1105), .B1(n4052), .C0(n891), 
        .C1(n4053), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[145]) );
  XOR2X1 U3301 ( .A(n4054), .B(n4055), .Y(n4053) );
  XOR2X1 U3302 ( .A(n4015), .B(n4048), .Y(n4055) );
  XNOR2X1 U3303 ( .A(n4056), .B(n3277), .Y(n4015) );
  XOR2X1 U3304 ( .A(n1392), .B(n1456), .Y(n3277) );
  CLKNAND2X2 U3305 ( .A(n1328), .B(n426), .Y(n4056) );
  AOI21X1 U3306 ( .A0(n924), .A1(n1386), .B0(n867), .Y(n4052) );
  AOI21X1 U3307 ( .A0(n1105), .A1(n931), .B0(n953), .Y(n4051) );
  OAI222X1 U3308 ( .A0(n1385), .A1(n4057), .B0(n1109), .B1(n4058), .C0(n891), 
        .C1(n4059), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[144]) );
  XOR2X1 U3309 ( .A(n4060), .B(n4061), .Y(n4059) );
  XOR2X1 U3310 ( .A(n4021), .B(n4054), .Y(n4061) );
  XNOR2X1 U3311 ( .A(n4062), .B(n3289), .Y(n4021) );
  XOR2X1 U3312 ( .A(n1391), .B(n1455), .Y(n3289) );
  CLKNAND2X2 U3313 ( .A(n1327), .B(n427), .Y(n4062) );
  AOI21X1 U3314 ( .A0(n927), .A1(n1385), .B0(n867), .Y(n4058) );
  AOI21X1 U3315 ( .A0(n1109), .A1(n931), .B0(n953), .Y(n4057) );
  OAI222X1 U3316 ( .A0(n1384), .A1(n4063), .B0(n1113), .B1(n4064), .C0(n891), 
        .C1(n4065), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[143]) );
  XOR2X1 U3317 ( .A(n4066), .B(n4067), .Y(n4065) );
  XOR2X1 U3318 ( .A(n4030), .B(n4060), .Y(n4067) );
  XNOR2X1 U3319 ( .A(n4068), .B(n3301), .Y(n4030) );
  XOR2X1 U3320 ( .A(n1390), .B(n1454), .Y(n3301) );
  CLKNAND2X2 U3321 ( .A(n1326), .B(n428), .Y(n4068) );
  AOI21X1 U3322 ( .A0(n927), .A1(n1384), .B0(n867), .Y(n4064) );
  AOI21X1 U3323 ( .A0(n1113), .A1(n931), .B0(n953), .Y(n4063) );
  OAI222X1 U3324 ( .A0(n1383), .A1(n4069), .B0(n1117), .B1(n4070), .C0(n891), 
        .C1(n4071), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[142]) );
  XOR2X1 U3325 ( .A(n4072), .B(n4073), .Y(n4071) );
  XOR2X1 U3326 ( .A(n4036), .B(n4066), .Y(n4073) );
  XNOR2X1 U3327 ( .A(n4074), .B(n3319), .Y(n4036) );
  XOR2X1 U3328 ( .A(n1389), .B(n1453), .Y(n3319) );
  CLKNAND2X2 U3329 ( .A(n1325), .B(n339), .Y(n4074) );
  AOI21X1 U3330 ( .A0(n925), .A1(n1383), .B0(n867), .Y(n4070) );
  AOI21X1 U3331 ( .A0(n1117), .A1(n930), .B0(n953), .Y(n4069) );
  OAI222X1 U3332 ( .A0(n1382), .A1(n4075), .B0(n1121), .B1(n4076), .C0(n891), 
        .C1(n4077), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[141]) );
  XOR2X1 U3333 ( .A(n4078), .B(n4079), .Y(n4077) );
  XOR2X1 U3334 ( .A(n4042), .B(n4072), .Y(n4079) );
  XNOR2X1 U3335 ( .A(n4080), .B(n3337), .Y(n4042) );
  XOR2X1 U3336 ( .A(n1388), .B(n1452), .Y(n3337) );
  CLKNAND2X2 U3337 ( .A(n1324), .B(n340), .Y(n4080) );
  AOI21X1 U3338 ( .A0(n927), .A1(n1382), .B0(n867), .Y(n4076) );
  AOI21X1 U3339 ( .A0(n1121), .A1(n930), .B0(n953), .Y(n4075) );
  OAI222X1 U3340 ( .A0(n1381), .A1(n4081), .B0(n1125), .B1(n4082), .C0(n891), 
        .C1(n4083), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[140]) );
  XOR2X1 U3341 ( .A(n4084), .B(n4085), .Y(n4083) );
  XOR2X1 U3342 ( .A(n4048), .B(n4078), .Y(n4085) );
  XNOR2X1 U3343 ( .A(n4086), .B(n3357), .Y(n4048) );
  XOR2X1 U3344 ( .A(n1387), .B(n1451), .Y(n3357) );
  CLKNAND2X2 U3345 ( .A(n1323), .B(n429), .Y(n4086) );
  AOI21X1 U3346 ( .A0(n924), .A1(n1381), .B0(n868), .Y(n4082) );
  AOI21X1 U3347 ( .A0(n1125), .A1(n930), .B0(n952), .Y(n4081) );
  OAI222X1 U3348 ( .A0(n878), .A1(n4087), .B0(n4088), .B1(n907), .C0(
        Inst_AEAD_u_input_n309), .C1(n856), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[13]) );
  XNOR2X1 U3349 ( .A(n2219), .B(n4089), .Y(n4088) );
  XOR2X1 U3350 ( .A(n2057), .B(n2164), .Y(n4089) );
  MXI2X1 U3351 ( .A(n2562), .B(n3429), .S0(n1487), .Y(n2164) );
  XNOR2X1 U3352 ( .A(n1359), .B(n1551), .Y(n2562) );
  MXI2X1 U3353 ( .A(n2709), .B(n4090), .S0(n1446), .Y(n2057) );
  XNOR2X1 U3354 ( .A(n1318), .B(n1510), .Y(n2709) );
  MXI2X1 U3355 ( .A(n2889), .B(n2081), .S0(n1453), .Y(n2219) );
  XNOR2X1 U3356 ( .A(n339), .B(n443), .Y(n2081) );
  XOR2X1 U3357 ( .A(n1325), .B(n1517), .Y(n2889) );
  OAI222X1 U3358 ( .A0(n1380), .A1(n4091), .B0(n1129), .B1(n4092), .C0(n891), 
        .C1(n4093), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[139]) );
  XNOR2X1 U3359 ( .A(n4094), .B(n4095), .Y(n4093) );
  XOR2X1 U3360 ( .A(n4054), .B(n4084), .Y(n4095) );
  XNOR2X1 U3361 ( .A(n4096), .B(n3381), .Y(n4054) );
  XOR2X1 U3362 ( .A(n1386), .B(n1450), .Y(n3381) );
  CLKNAND2X2 U3363 ( .A(n1322), .B(n430), .Y(n4096) );
  AOI21X1 U3364 ( .A0(n925), .A1(n1380), .B0(n868), .Y(n4092) );
  AOI21X1 U3365 ( .A0(n1129), .A1(n929), .B0(n952), .Y(n4091) );
  OAI222X1 U3366 ( .A0(n1379), .A1(n4097), .B0(n1133), .B1(n4098), .C0(n892), 
        .C1(n4099), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[138]) );
  XOR2X1 U3367 ( .A(n4100), .B(n4101), .Y(n4099) );
  XNOR2X1 U3368 ( .A(n4060), .B(n4094), .Y(n4101) );
  CLKINVX1 U3369 ( .A(n4102), .Y(n4094) );
  XNOR2X1 U3370 ( .A(n4103), .B(n4104), .Y(n4060) );
  CLKNAND2X2 U3371 ( .A(n1321), .B(n406), .Y(n4103) );
  AOI21X1 U3372 ( .A0(n926), .A1(n1379), .B0(n868), .Y(n4098) );
  AOI21X1 U3373 ( .A0(n1133), .A1(n931), .B0(n952), .Y(n4097) );
  OAI222X1 U3374 ( .A0(n1378), .A1(n4105), .B0(n1137), .B1(n4106), .C0(n892), 
        .C1(n4107), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[137]) );
  XOR2X1 U3375 ( .A(n4108), .B(n4109), .Y(n4107) );
  XOR2X1 U3376 ( .A(n4066), .B(n4100), .Y(n4109) );
  XNOR2X1 U3377 ( .A(n4110), .B(n4111), .Y(n4066) );
  CLKNAND2X2 U3378 ( .A(n1320), .B(n407), .Y(n4110) );
  AOI21X1 U3379 ( .A0(n926), .A1(n1378), .B0(n868), .Y(n4106) );
  AOI21X1 U3380 ( .A0(n1137), .A1(n930), .B0(n952), .Y(n4105) );
  OAI222X1 U3381 ( .A0(n1377), .A1(n4112), .B0(n1141), .B1(n4113), .C0(n892), 
        .C1(n4114), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[136]) );
  XNOR2X1 U3382 ( .A(n4115), .B(n4116), .Y(n4114) );
  XOR2X1 U3383 ( .A(n4072), .B(n4108), .Y(n4116) );
  XNOR2X1 U3384 ( .A(n4117), .B(n4118), .Y(n4072) );
  CLKNAND2X2 U3385 ( .A(n1319), .B(n408), .Y(n4117) );
  AOI21X1 U3386 ( .A0(n925), .A1(n1377), .B0(n868), .Y(n4113) );
  AOI21X1 U3387 ( .A0(n1141), .A1(n929), .B0(n952), .Y(n4112) );
  OAI222X1 U3388 ( .A0(n1376), .A1(n4119), .B0(n1145), .B1(n4120), .C0(n889), 
        .C1(n4121), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[135]) );
  XNOR2X1 U3389 ( .A(n4122), .B(n4123), .Y(n4121) );
  XNOR2X1 U3390 ( .A(n4124), .B(n4078), .Y(n4123) );
  XNOR2X1 U3391 ( .A(n4125), .B(n4126), .Y(n4078) );
  CLKNAND2X2 U3392 ( .A(n1318), .B(n431), .Y(n4125) );
  AOI21X1 U3393 ( .A0(n926), .A1(n1376), .B0(n868), .Y(n4120) );
  AOI21X1 U3394 ( .A0(n1145), .A1(n929), .B0(n952), .Y(n4119) );
  OAI222X1 U3395 ( .A0(n1375), .A1(n4127), .B0(n1149), .B1(n4128), .C0(n892), 
        .C1(n4129), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[134]) );
  XNOR2X1 U3396 ( .A(n4130), .B(n4131), .Y(n4129) );
  XNOR2X1 U3397 ( .A(n4122), .B(n4084), .Y(n4131) );
  XNOR2X1 U3398 ( .A(n4132), .B(n4133), .Y(n4084) );
  CLKNAND2X2 U3399 ( .A(n1317), .B(n432), .Y(n4132) );
  AOI21X1 U3400 ( .A0(n926), .A1(n1375), .B0(n868), .Y(n4128) );
  AOI21X1 U3401 ( .A0(n1149), .A1(n928), .B0(n952), .Y(n4127) );
  OAI222X1 U3402 ( .A0(n1374), .A1(n4134), .B0(n1153), .B1(n4135), .C0(n892), 
        .C1(n4136), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[133]) );
  XOR2X1 U3403 ( .A(n4130), .B(n4137), .Y(n4136) );
  XNOR2X1 U3404 ( .A(n3742), .B(n4102), .Y(n4137) );
  XOR2X1 U3405 ( .A(n4138), .B(n3494), .Y(n4102) );
  CLKNAND2X2 U3406 ( .A(n1316), .B(n433), .Y(n4138) );
  AOI21X1 U3407 ( .A0(n924), .A1(n1374), .B0(n868), .Y(n4135) );
  AOI21X1 U3408 ( .A0(n1153), .A1(n928), .B0(n952), .Y(n4134) );
  OAI222X1 U3409 ( .A0(n1373), .A1(n4139), .B0(n1157), .B1(n4140), .C0(n892), 
        .C1(n4141), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[132]) );
  XOR2X1 U3410 ( .A(n4100), .B(n4142), .Y(n4141) );
  XOR2X1 U3411 ( .A(n3742), .B(n3749), .Y(n4142) );
  XOR2X1 U3412 ( .A(n3621), .B(n4143), .Y(n3742) );
  NOR2X1 U3413 ( .A(n1247), .B(n436), .Y(n4143) );
  XNOR2X1 U3414 ( .A(n4144), .B(n4145), .Y(n4100) );
  CLKNAND2X2 U3415 ( .A(n1315), .B(n434), .Y(n4144) );
  AOI21X1 U3416 ( .A0(n925), .A1(n1373), .B0(n868), .Y(n4140) );
  AOI21X1 U3417 ( .A0(n1157), .A1(n929), .B0(n952), .Y(n4139) );
  OAI222X1 U3418 ( .A0(n1372), .A1(n4146), .B0(n1161), .B1(n4147), .C0(n892), 
        .C1(n4148), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[131]) );
  XOR2X1 U3419 ( .A(n4108), .B(n4149), .Y(n4148) );
  XOR2X1 U3420 ( .A(n3749), .B(n3758), .Y(n4149) );
  XOR2X1 U3421 ( .A(n3640), .B(n4150), .Y(n3749) );
  NOR2X1 U3422 ( .A(n1246), .B(n437), .Y(n4150) );
  XNOR2X1 U3423 ( .A(n4151), .B(n4152), .Y(n4108) );
  CLKNAND2X2 U3424 ( .A(n1314), .B(n409), .Y(n4151) );
  AOI21X1 U3425 ( .A0(n925), .A1(n1372), .B0(n868), .Y(n4147) );
  AOI21X1 U3426 ( .A0(n1161), .A1(n928), .B0(n952), .Y(n4146) );
  OAI222X1 U3427 ( .A0(n1371), .A1(n4153), .B0(n1165), .B1(n4154), .C0(n892), 
        .C1(n4155), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[130]) );
  XNOR2X1 U3428 ( .A(n4115), .B(n4156), .Y(n4155) );
  XOR2X1 U3429 ( .A(n3758), .B(n3764), .Y(n4156) );
  XOR2X1 U3430 ( .A(n3659), .B(n4157), .Y(n3758) );
  NOR2X1 U3431 ( .A(n1245), .B(n438), .Y(n4157) );
  CLKINVX1 U3432 ( .A(n4124), .Y(n4115) );
  XOR2X1 U3433 ( .A(n4158), .B(n3548), .Y(n4124) );
  CLKNAND2X2 U3434 ( .A(n1313), .B(n410), .Y(n4158) );
  AOI21X1 U3435 ( .A0(n924), .A1(n1371), .B0(n868), .Y(n4154) );
  AOI21X1 U3436 ( .A0(n1165), .A1(n928), .B0(n952), .Y(n4153) );
  OAI222X1 U3437 ( .A0(n877), .A1(n4159), .B0(n903), .B1(n4160), .C0(
        Inst_AEAD_u_input_n310), .C1(n854), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[12]) );
  XNOR2X1 U3438 ( .A(n2226), .B(n4161), .Y(n4160) );
  XOR2X1 U3439 ( .A(n2169), .B(n2132), .Y(n4161) );
  MXI2X1 U3440 ( .A(n2721), .B(n4162), .S0(n1445), .Y(n2132) );
  XNOR2X1 U3441 ( .A(n1317), .B(n1509), .Y(n2721) );
  MXI2X1 U3442 ( .A(n2570), .B(n3449), .S0(n1486), .Y(n2169) );
  XOR2X1 U3443 ( .A(n1358), .B(n347), .Y(n2570) );
  MXI2X1 U3444 ( .A(n2908), .B(n2089), .S0(n1452), .Y(n2226) );
  XNOR2X1 U3445 ( .A(n340), .B(n444), .Y(n2089) );
  XOR2X1 U3446 ( .A(n1324), .B(n1516), .Y(n2908) );
  OAI222X1 U3447 ( .A0(n1370), .A1(n4163), .B0(n1169), .B1(n4164), .C0(n892), 
        .C1(n4165), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[129]) );
  XOR2X1 U3448 ( .A(n4122), .B(n4166), .Y(n4165) );
  XOR2X1 U3449 ( .A(n3764), .B(n3770), .Y(n4166) );
  XOR2X1 U3450 ( .A(n3685), .B(n4167), .Y(n3764) );
  NOR2X1 U3451 ( .A(n1244), .B(n439), .Y(n4167) );
  XNOR2X1 U3452 ( .A(n3583), .B(n4168), .Y(n4122) );
  NOR2X1 U3453 ( .A(n1249), .B(n441), .Y(n4168) );
  AOI21X1 U3454 ( .A0(n924), .A1(n1370), .B0(n868), .Y(n4164) );
  AOI21X1 U3455 ( .A0(n1169), .A1(n929), .B0(n952), .Y(n4163) );
  OAI222X1 U3456 ( .A0(n1369), .A1(n4169), .B0(n1173), .B1(n4170), .C0(n887), 
        .C1(n4171), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[128]) );
  XOR2X1 U3457 ( .A(n4130), .B(n4172), .Y(n4171) );
  XOR2X1 U3458 ( .A(n3744), .B(n3770), .Y(n4172) );
  XOR2X1 U3459 ( .A(n3710), .B(n4173), .Y(n3770) );
  NOR2X1 U3460 ( .A(n1243), .B(n440), .Y(n4173) );
  XOR2X1 U3461 ( .A(n3734), .B(n4174), .Y(n3744) );
  AND2X1 U3462 ( .A(n1241), .B(n378), .Y(n4174) );
  XNOR2X1 U3463 ( .A(n3602), .B(n4175), .Y(n4130) );
  NOR2X1 U3464 ( .A(n1248), .B(n435), .Y(n4175) );
  AOI21X1 U3465 ( .A0(n924), .A1(n1369), .B0(n868), .Y(n4170) );
  AOI21X1 U3466 ( .A0(n1173), .A1(n927), .B0(n952), .Y(n4169) );
  NOR2X1 U3467 ( .A(n879), .B(n927), .Y(n2923) );
  OAI222X1 U3468 ( .A0(n878), .A1(n4176), .B0(n903), .B1(n4177), .C0(n1177), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[127]) );
  XNOR2X1 U3469 ( .A(n4178), .B(n4179), .Y(n4177) );
  XOR2X1 U3470 ( .A(n1969), .B(n2025), .Y(n4179) );
  XNOR2X1 U3471 ( .A(n3396), .B(n4180), .Y(n1969) );
  NOR2X1 U3472 ( .A(n348), .B(n3401), .Y(n4180) );
  XOR2X1 U3473 ( .A(n1258), .B(n1321), .Y(n3401) );
  CLKINVX1 U3474 ( .A(n4104), .Y(n3396) );
  XOR2X1 U3475 ( .A(n1385), .B(n1449), .Y(n4104) );
  OAI222X1 U3476 ( .A0(n878), .A1(n4181), .B0(n903), .B1(n4182), .C0(n1178), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[126]) );
  XNOR2X1 U3477 ( .A(n4183), .B(n4184), .Y(n4182) );
  XOR2X1 U3478 ( .A(n1983), .B(n2032), .Y(n4184) );
  XNOR2X1 U3479 ( .A(n3416), .B(n4185), .Y(n1983) );
  NOR2X1 U3480 ( .A(n349), .B(n3421), .Y(n4185) );
  XOR2X1 U3481 ( .A(n1257), .B(n1320), .Y(n3421) );
  CLKINVX1 U3482 ( .A(n4111), .Y(n3416) );
  XOR2X1 U3483 ( .A(n1384), .B(n1448), .Y(n4111) );
  OAI222X1 U3484 ( .A0(n878), .A1(n4186), .B0(n904), .B1(n4187), .C0(n1179), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[125]) );
  XNOR2X1 U3485 ( .A(n4188), .B(n4189), .Y(n4187) );
  XNOR2X1 U3486 ( .A(n2044), .B(n1990), .Y(n4189) );
  XNOR2X1 U3487 ( .A(n3436), .B(n4190), .Y(n1990) );
  NOR2X1 U3488 ( .A(n3441), .B(n371), .Y(n4190) );
  XOR2X1 U3489 ( .A(n1256), .B(n1319), .Y(n3441) );
  CLKINVX1 U3490 ( .A(n4118), .Y(n3436) );
  XOR2X1 U3491 ( .A(n1383), .B(n1447), .Y(n4118) );
  OAI222X1 U3492 ( .A0(n878), .A1(n4191), .B0(n903), .B1(n4192), .C0(n1180), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[124]) );
  XNOR2X1 U3493 ( .A(n4193), .B(n4194), .Y(n4192) );
  XNOR2X1 U3494 ( .A(n2052), .B(n1997), .Y(n4194) );
  XNOR2X1 U3495 ( .A(n3456), .B(n4195), .Y(n1997) );
  AND2X1 U3496 ( .A(n1510), .B(n2712), .Y(n4195) );
  CLKINVX1 U3497 ( .A(n4090), .Y(n2712) );
  XNOR2X1 U3498 ( .A(n1255), .B(n460), .Y(n4090) );
  CLKINVX1 U3499 ( .A(n4126), .Y(n3456) );
  XOR2X1 U3500 ( .A(n1382), .B(n1446), .Y(n4126) );
  OAI222X1 U3501 ( .A0(n878), .A1(n4196), .B0(n904), .B1(n4197), .C0(n1181), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[123]) );
  XNOR2X1 U3502 ( .A(n4198), .B(n4199), .Y(n4197) );
  XNOR2X1 U3503 ( .A(n2066), .B(n2004), .Y(n4199) );
  XNOR2X1 U3504 ( .A(n3475), .B(n4200), .Y(n2004) );
  AND2X1 U3505 ( .A(n1509), .B(n2724), .Y(n4200) );
  CLKINVX1 U3506 ( .A(n4162), .Y(n2724) );
  XNOR2X1 U3507 ( .A(n1254), .B(n461), .Y(n4162) );
  CLKINVX1 U3508 ( .A(n4133), .Y(n3475) );
  XOR2X1 U3509 ( .A(n1381), .B(n1445), .Y(n4133) );
  OAI222X1 U3510 ( .A0(n878), .A1(n4201), .B0(n903), .B1(n4202), .C0(n1182), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[122]) );
  XNOR2X1 U3511 ( .A(n4203), .B(n4204), .Y(n4202) );
  XNOR2X1 U3512 ( .A(n2074), .B(n2011), .Y(n4204) );
  XNOR2X1 U3513 ( .A(n3494), .B(n4205), .Y(n2011) );
  AND2X1 U3514 ( .A(n1508), .B(n2735), .Y(n4205) );
  CLKINVX1 U3515 ( .A(n4206), .Y(n2735) );
  XNOR2X1 U3516 ( .A(n1380), .B(n1444), .Y(n3494) );
  OAI222X1 U3517 ( .A0(n878), .A1(n4207), .B0(n904), .B1(n4208), .C0(n1183), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[121]) );
  XNOR2X1 U3518 ( .A(n4209), .B(n4210), .Y(n4208) );
  XNOR2X1 U3519 ( .A(n2082), .B(n2018), .Y(n4210) );
  XNOR2X1 U3520 ( .A(n3512), .B(n4211), .Y(n2018) );
  AND2X1 U3521 ( .A(n1507), .B(n2746), .Y(n4211) );
  CLKINVX1 U3522 ( .A(n4212), .Y(n2746) );
  CLKINVX1 U3523 ( .A(n4145), .Y(n3512) );
  XOR2X1 U3524 ( .A(n1379), .B(n1443), .Y(n4145) );
  OAI222X1 U3525 ( .A0(n878), .A1(n4213), .B0(n903), .B1(n4214), .C0(n1184), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[120]) );
  XNOR2X1 U3526 ( .A(n4215), .B(n4216), .Y(n4214) );
  XNOR2X1 U3527 ( .A(n2090), .B(n2025), .Y(n4216) );
  XNOR2X1 U3528 ( .A(n3530), .B(n4217), .Y(n2025) );
  NOR2X1 U3529 ( .A(n2417), .B(n372), .Y(n4217) );
  XOR2X1 U3530 ( .A(n1251), .B(n1314), .Y(n2417) );
  CLKINVX1 U3531 ( .A(n4152), .Y(n3530) );
  XOR2X1 U3532 ( .A(n1378), .B(n1442), .Y(n4152) );
  OAI222X1 U3533 ( .A0(n878), .A1(n4218), .B0(n904), .B1(n4219), .C0(
        Inst_AEAD_u_input_n311), .C1(n856), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[11]) );
  XOR2X1 U3534 ( .A(n2234), .B(n4220), .Y(n4219) );
  XOR2X1 U3535 ( .A(n2188), .B(n2175), .Y(n4220) );
  MXI2X1 U3536 ( .A(n2580), .B(n3468), .S0(n1485), .Y(n2175) );
  XOR2X1 U3537 ( .A(n1357), .B(n359), .Y(n2580) );
  MXI2X1 U3538 ( .A(n2732), .B(n4206), .S0(n1444), .Y(n2188) );
  XNOR2X1 U3539 ( .A(n1253), .B(n462), .Y(n4206) );
  XNOR2X1 U3540 ( .A(n1316), .B(n1508), .Y(n2732) );
  MXI2X1 U3541 ( .A(n2639), .B(n3356), .S0(n1451), .Y(n2234) );
  XNOR2X1 U3542 ( .A(n1260), .B(n463), .Y(n3356) );
  XNOR2X1 U3543 ( .A(n1323), .B(n1515), .Y(n2639) );
  OAI222X1 U3544 ( .A0(n878), .A1(n4221), .B0(n902), .B1(n4222), .C0(n1185), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[119]) );
  XNOR2X1 U3545 ( .A(n4223), .B(n4224), .Y(n4222) );
  XNOR2X1 U3546 ( .A(n2098), .B(n2032), .Y(n4224) );
  XNOR2X1 U3547 ( .A(n3548), .B(n4225), .Y(n2032) );
  NOR2X1 U3548 ( .A(n3553), .B(n373), .Y(n4225) );
  XOR2X1 U3549 ( .A(n1250), .B(n1313), .Y(n3553) );
  XNOR2X1 U3550 ( .A(n1377), .B(n1441), .Y(n3548) );
  OAI222X1 U3551 ( .A0(n878), .A1(n4226), .B0(n904), .B1(n4227), .C0(n1186), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[118]) );
  XOR2X1 U3552 ( .A(n4228), .B(n4229), .Y(n4227) );
  XNOR2X1 U3553 ( .A(n2044), .B(n2101), .Y(n4229) );
  CLKINVX1 U3554 ( .A(n4230), .Y(n2101) );
  XNOR2X1 U3555 ( .A(n3583), .B(n4231), .Y(n2044) );
  NOR2X1 U3556 ( .A(n350), .B(n4232), .Y(n4231) );
  XNOR2X1 U3557 ( .A(n1440), .B(n2785), .Y(n3583) );
  XOR2X1 U3558 ( .A(Inst_AEAD_u_cc_u_cc_dp_rc_7_), .B(n1376), .Y(n2785) );
  OAI222X1 U3559 ( .A0(n878), .A1(n4233), .B0(n904), .B1(n4234), .C0(n1187), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[117]) );
  XOR2X1 U3560 ( .A(n4235), .B(n4236), .Y(n4234) );
  XNOR2X1 U3561 ( .A(n2052), .B(n4178), .Y(n4236) );
  XNOR2X1 U3562 ( .A(n3602), .B(n4237), .Y(n2052) );
  AND2X1 U3563 ( .A(n1503), .B(n2423), .Y(n4237) );
  XOR2X1 U3564 ( .A(n1248), .B(n435), .Y(n2423) );
  XNOR2X1 U3565 ( .A(n1439), .B(n2801), .Y(n3602) );
  XNOR2X1 U3566 ( .A(n377), .B(n1375), .Y(n2801) );
  OAI222X1 U3567 ( .A0(n878), .A1(n4238), .B0(n903), .B1(n4239), .C0(n1188), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[116]) );
  XNOR2X1 U3568 ( .A(n4240), .B(n4241), .Y(n4239) );
  XNOR2X1 U3569 ( .A(n2066), .B(n1867), .Y(n4241) );
  XNOR2X1 U3570 ( .A(n3621), .B(n4242), .Y(n2066) );
  AND2X1 U3571 ( .A(n1502), .B(n2491), .Y(n4242) );
  XOR2X1 U3572 ( .A(n1247), .B(n436), .Y(n2491) );
  XNOR2X1 U3573 ( .A(n1438), .B(n2817), .Y(n3621) );
  XOR2X1 U3574 ( .A(n1374), .B(Inst_AEAD_u_cc_u_cc_dp_rc_5_), .Y(n2817) );
  OAI222X1 U3575 ( .A0(n878), .A1(n4243), .B0(n904), .B1(n4244), .C0(n1189), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[115]) );
  XNOR2X1 U3576 ( .A(n4188), .B(n4245), .Y(n4244) );
  XNOR2X1 U3577 ( .A(n2074), .B(n1873), .Y(n4245) );
  XNOR2X1 U3578 ( .A(n3640), .B(n4246), .Y(n2074) );
  AND2X1 U3579 ( .A(n1501), .B(n2590), .Y(n4246) );
  XOR2X1 U3580 ( .A(n1246), .B(n437), .Y(n2590) );
  XNOR2X1 U3581 ( .A(n1437), .B(n2833), .Y(n3640) );
  XOR2X1 U3582 ( .A(n1373), .B(Inst_AEAD_u_cc_u_cc_dp_rc_4_), .Y(n2833) );
  OAI222X1 U3583 ( .A0(n878), .A1(n4247), .B0(n902), .B1(n4248), .C0(n1190), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[114]) );
  XNOR2X1 U3584 ( .A(n4193), .B(n4249), .Y(n4248) );
  XNOR2X1 U3585 ( .A(n2082), .B(n1879), .Y(n4249) );
  XNOR2X1 U3586 ( .A(n3659), .B(n4250), .Y(n2082) );
  AND2X1 U3587 ( .A(n1500), .B(n2699), .Y(n4250) );
  XOR2X1 U3588 ( .A(n1245), .B(n438), .Y(n2699) );
  XNOR2X1 U3589 ( .A(n1436), .B(n2856), .Y(n3659) );
  XOR2X1 U3590 ( .A(Inst_AEAD_u_cc_u_cc_dp_rc_3_), .B(n1372), .Y(n2856) );
  OAI222X1 U3591 ( .A0(n878), .A1(n4251), .B0(n904), .B1(n4252), .C0(n1191), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[113]) );
  XNOR2X1 U3592 ( .A(n4198), .B(n4253), .Y(n4252) );
  XNOR2X1 U3593 ( .A(n2090), .B(n1885), .Y(n4253) );
  XNOR2X1 U3594 ( .A(n3685), .B(n4254), .Y(n2090) );
  AND2X1 U3595 ( .A(n1499), .B(n2849), .Y(n4254) );
  XOR2X1 U3596 ( .A(n1244), .B(n439), .Y(n2849) );
  XNOR2X1 U3597 ( .A(n1435), .B(n2871), .Y(n3685) );
  XOR2X1 U3598 ( .A(n1371), .B(Inst_AEAD_u_cc_u_cc_dp_rc_2_), .Y(n2871) );
  OAI222X1 U3599 ( .A0(n879), .A1(n4255), .B0(n903), .B1(n4256), .C0(n1192), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[112]) );
  XNOR2X1 U3600 ( .A(n4203), .B(n4257), .Y(n4256) );
  XNOR2X1 U3601 ( .A(n2098), .B(n1891), .Y(n4257) );
  XNOR2X1 U3602 ( .A(n3710), .B(n4258), .Y(n2098) );
  AND2X1 U3603 ( .A(n1498), .B(n2886), .Y(n4258) );
  XOR2X1 U3604 ( .A(n1243), .B(n440), .Y(n2886) );
  XNOR2X1 U3605 ( .A(n1434), .B(n2888), .Y(n3710) );
  XOR2X1 U3606 ( .A(n1370), .B(Inst_AEAD_u_cc_u_cc_dp_rc_1_), .Y(n2888) );
  OAI222X1 U3607 ( .A0(n878), .A1(n4259), .B0(n902), .B1(n4260), .C0(n1193), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[111]) );
  XNOR2X1 U3608 ( .A(n4209), .B(n4261), .Y(n4260) );
  XNOR2X1 U3609 ( .A(n4230), .B(n1897), .Y(n4261) );
  XNOR2X1 U3610 ( .A(n3734), .B(n4262), .Y(n4230) );
  AND2X1 U3611 ( .A(n1497), .B(n2905), .Y(n4262) );
  XNOR2X1 U3612 ( .A(n1433), .B(n2907), .Y(n3734) );
  XOR2X1 U3613 ( .A(n1369), .B(Inst_AEAD_u_cc_u_cc_dp_rc_0_), .Y(n2907) );
  OAI222X1 U3614 ( .A0(n878), .A1(n4263), .B0(n903), .B1(n4264), .C0(n1194), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[110]) );
  XOR2X1 U3615 ( .A(n4215), .B(n4265), .Y(n4264) );
  XNOR2X1 U3616 ( .A(n1903), .B(n4178), .Y(n4265) );
  XOR2X1 U3617 ( .A(n3678), .B(n4266), .Y(n4178) );
  NOR2BX1 U3618 ( .AN(n1560), .B(n3089), .Y(n4266) );
  XOR2X1 U3619 ( .A(n1305), .B(n1368), .Y(n3089) );
  XNOR2X1 U3620 ( .A(n1432), .B(n1496), .Y(n3678) );
  OAI222X1 U3621 ( .A0(n879), .A1(n4267), .B0(n4268), .B1(n906), .C0(
        Inst_AEAD_u_input_n312), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[10]) );
  XOR2X1 U3622 ( .A(n4269), .B(n2246), .Y(n4268) );
  MXI2X1 U3623 ( .A(n2743), .B(n4212), .S0(n1443), .Y(n2246) );
  XNOR2X1 U3624 ( .A(n1252), .B(n464), .Y(n4212) );
  XNOR2X1 U3625 ( .A(n1315), .B(n1507), .Y(n2743) );
  XOR2X1 U3626 ( .A(n2239), .B(n2180), .Y(n4269) );
  MXI2X1 U3627 ( .A(n2599), .B(n3487), .S0(n1484), .Y(n2180) );
  XOR2X1 U3628 ( .A(n1356), .B(n361), .Y(n2599) );
  MXI2X1 U3629 ( .A(n2650), .B(n3380), .S0(n1450), .Y(n2239) );
  XNOR2X1 U3630 ( .A(n1259), .B(n465), .Y(n3380) );
  XNOR2X1 U3631 ( .A(n1322), .B(n1514), .Y(n2650) );
  OAI222X1 U3632 ( .A0(n879), .A1(n4270), .B0(n902), .B1(n4271), .C0(n1195), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[109]) );
  XOR2X1 U3633 ( .A(n4223), .B(n4272), .Y(n4271) );
  XNOR2X1 U3634 ( .A(n1866), .B(n4183), .Y(n4272) );
  CLKINVX1 U3635 ( .A(n4240), .Y(n4183) );
  XOR2X1 U3636 ( .A(n3790), .B(n4273), .Y(n4240) );
  NOR2X1 U3637 ( .A(n3214), .B(n354), .Y(n4273) );
  XOR2X1 U3638 ( .A(n1304), .B(n1367), .Y(n3214) );
  XOR2X1 U3639 ( .A(n1431), .B(n1495), .Y(n3790) );
  XNOR2X1 U3640 ( .A(n3595), .B(n4274), .Y(n1866) );
  NOR2X1 U3641 ( .A(n2256), .B(n355), .Y(n4274) );
  XOR2X1 U3642 ( .A(n1287), .B(n1350), .Y(n2256) );
  CLKINVX1 U3643 ( .A(n3909), .Y(n3595) );
  XOR2X1 U3644 ( .A(n1414), .B(n1478), .Y(n3909) );
  OAI222X1 U3645 ( .A0(n879), .A1(n4275), .B0(n904), .B1(n4276), .C0(n1196), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[108]) );
  XOR2X1 U3646 ( .A(n4228), .B(n4277), .Y(n4276) );
  XOR2X1 U3647 ( .A(n1872), .B(n4188), .Y(n4277) );
  XOR2X1 U3648 ( .A(n3797), .B(n4278), .Y(n4188) );
  NOR2X1 U3649 ( .A(n3369), .B(n356), .Y(n4278) );
  XOR2X1 U3650 ( .A(n1303), .B(n1366), .Y(n3369) );
  XOR2X1 U3651 ( .A(n1430), .B(n1494), .Y(n3797) );
  XNOR2X1 U3652 ( .A(n3614), .B(n4279), .Y(n1872) );
  NOR2X1 U3653 ( .A(n2261), .B(n357), .Y(n4279) );
  XOR2X1 U3654 ( .A(n1286), .B(n1349), .Y(n2261) );
  CLKINVX1 U3655 ( .A(n3916), .Y(n3614) );
  XOR2X1 U3656 ( .A(n1413), .B(n1477), .Y(n3916) );
  OAI222X1 U3657 ( .A0(n879), .A1(n4280), .B0(n904), .B1(n4281), .C0(n1197), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[107]) );
  XOR2X1 U3658 ( .A(n4235), .B(n4282), .Y(n4281) );
  XOR2X1 U3659 ( .A(n1878), .B(n4193), .Y(n4282) );
  XOR2X1 U3660 ( .A(n3804), .B(n4283), .Y(n4193) );
  NOR2X1 U3661 ( .A(n3309), .B(n358), .Y(n4283) );
  XOR2X1 U3662 ( .A(n1302), .B(n1365), .Y(n3309) );
  XOR2X1 U3663 ( .A(n1429), .B(n1493), .Y(n3804) );
  XNOR2X1 U3664 ( .A(n3633), .B(n4284), .Y(n1878) );
  NOR2X1 U3665 ( .A(n2415), .B(n379), .Y(n4284) );
  XOR2X1 U3666 ( .A(n1285), .B(n1348), .Y(n2415) );
  CLKINVX1 U3667 ( .A(n3923), .Y(n3633) );
  XOR2X1 U3668 ( .A(n1412), .B(n1476), .Y(n3923) );
  OAI222X1 U3669 ( .A0(n879), .A1(n4285), .B0(n904), .B1(n4286), .C0(n1198), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[106]) );
  XOR2X1 U3670 ( .A(n4198), .B(n4287), .Y(n4286) );
  XOR2X1 U3671 ( .A(n1867), .B(n1884), .Y(n4287) );
  XNOR2X1 U3672 ( .A(n3652), .B(n4288), .Y(n1884) );
  NOR2X1 U3673 ( .A(n3564), .B(n380), .Y(n4288) );
  XOR2X1 U3674 ( .A(n1284), .B(n1347), .Y(n3564) );
  CLKINVX1 U3675 ( .A(n3930), .Y(n3652) );
  XOR2X1 U3676 ( .A(n1411), .B(n1475), .Y(n3930) );
  XNOR2X1 U3677 ( .A(n3463), .B(n4289), .Y(n1867) );
  NOR2X1 U3678 ( .A(n3468), .B(n359), .Y(n4289) );
  XOR2X1 U3679 ( .A(n1294), .B(n1357), .Y(n3468) );
  CLKINVX1 U3680 ( .A(n3857), .Y(n3463) );
  XOR2X1 U3681 ( .A(n1421), .B(n1485), .Y(n3857) );
  XOR2X1 U3682 ( .A(n3811), .B(n4290), .Y(n4198) );
  NOR2X1 U3683 ( .A(n3327), .B(n360), .Y(n4290) );
  XOR2X1 U3684 ( .A(n1301), .B(n1364), .Y(n3327) );
  XOR2X1 U3685 ( .A(n1428), .B(n1492), .Y(n3811) );
  OAI222X1 U3686 ( .A0(n879), .A1(n4291), .B0(n905), .B1(n4292), .C0(n1199), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[105]) );
  XOR2X1 U3687 ( .A(n4203), .B(n4293), .Y(n4292) );
  XOR2X1 U3688 ( .A(n1873), .B(n1890), .Y(n4293) );
  XNOR2X1 U3689 ( .A(n3670), .B(n4294), .Y(n1890) );
  NOR2X1 U3690 ( .A(n3675), .B(n370), .Y(n4294) );
  CLKINVX1 U3691 ( .A(n3937), .Y(n3670) );
  XOR2X1 U3692 ( .A(n1410), .B(n1474), .Y(n3937) );
  XNOR2X1 U3693 ( .A(n3482), .B(n4295), .Y(n1873) );
  NOR2X1 U3694 ( .A(n3487), .B(n361), .Y(n4295) );
  XOR2X1 U3695 ( .A(n1293), .B(n1356), .Y(n3487) );
  CLKINVX1 U3696 ( .A(n3864), .Y(n3482) );
  XOR2X1 U3697 ( .A(n1420), .B(n1484), .Y(n3864) );
  XNOR2X1 U3698 ( .A(n3340), .B(n4296), .Y(n4203) );
  NOR2X1 U3699 ( .A(n3345), .B(n362), .Y(n4296) );
  XOR2X1 U3700 ( .A(n1300), .B(n1363), .Y(n3345) );
  XNOR2X1 U3701 ( .A(n1427), .B(n1491), .Y(n3340) );
  OAI222X1 U3702 ( .A0(n879), .A1(n4297), .B0(n903), .B1(n4298), .C0(n1200), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[104]) );
  XOR2X1 U3703 ( .A(n4209), .B(n4299), .Y(n4298) );
  XOR2X1 U3704 ( .A(n1879), .B(n1896), .Y(n4299) );
  XNOR2X1 U3705 ( .A(n3696), .B(n4300), .Y(n1896) );
  NOR2X1 U3706 ( .A(n2275), .B(n363), .Y(n4300) );
  XOR2X1 U3707 ( .A(n1282), .B(n1345), .Y(n2275) );
  CLKINVX1 U3708 ( .A(n3944), .Y(n3696) );
  XOR2X1 U3709 ( .A(n1409), .B(n1473), .Y(n3944) );
  XNOR2X1 U3710 ( .A(n3501), .B(n4301), .Y(n1879) );
  NOR2X1 U3711 ( .A(n2222), .B(n364), .Y(n4301) );
  XOR2X1 U3712 ( .A(n1292), .B(n1355), .Y(n2222) );
  CLKINVX1 U3713 ( .A(n3871), .Y(n3501) );
  XOR2X1 U3714 ( .A(n1419), .B(n1483), .Y(n3871) );
  XNOR2X1 U3715 ( .A(n3360), .B(n4302), .Y(n4209) );
  NOR2X1 U3716 ( .A(n344), .B(n3365), .Y(n4302) );
  XOR2X1 U3717 ( .A(n1299), .B(n1362), .Y(n3365) );
  XNOR2X1 U3718 ( .A(n1426), .B(n1490), .Y(n3360) );
  OAI222X1 U3719 ( .A0(n879), .A1(n4303), .B0(n905), .B1(n4304), .C0(n1201), 
        .C1(n855), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[103]) );
  XOR2X1 U3720 ( .A(n4215), .B(n4305), .Y(n4304) );
  XOR2X1 U3721 ( .A(n1885), .B(n1902), .Y(n4305) );
  XNOR2X1 U3722 ( .A(n3721), .B(n4306), .Y(n1902) );
  NOR2BX1 U3723 ( .AN(n2280), .B(n351), .Y(n4306) );
  XNOR2X1 U3724 ( .A(n1281), .B(n1344), .Y(n2280) );
  CLKINVX1 U3725 ( .A(n3951), .Y(n3721) );
  XOR2X1 U3726 ( .A(n1408), .B(n1472), .Y(n3951) );
  XNOR2X1 U3727 ( .A(n3519), .B(n4307), .Y(n1885) );
  NOR2X1 U3728 ( .A(n2229), .B(n365), .Y(n4307) );
  XOR2X1 U3729 ( .A(n1291), .B(n1354), .Y(n2229) );
  CLKINVX1 U3730 ( .A(n3878), .Y(n3519) );
  XOR2X1 U3731 ( .A(n1418), .B(n1482), .Y(n3878) );
  XNOR2X1 U3732 ( .A(n3384), .B(n4308), .Y(n4215) );
  NOR2X1 U3733 ( .A(n345), .B(n3389), .Y(n4308) );
  XOR2X1 U3734 ( .A(n1298), .B(n1361), .Y(n3389) );
  XNOR2X1 U3735 ( .A(n1425), .B(n1489), .Y(n3384) );
  OAI222X1 U3736 ( .A0(n879), .A1(n4309), .B0(n904), .B1(n4310), .C0(n1202), 
        .C1(n853), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[102]) );
  XOR2X1 U3737 ( .A(n4223), .B(n4311), .Y(n4310) );
  XOR2X1 U3738 ( .A(n1891), .B(n1906), .Y(n4311) );
  XNOR2X1 U3739 ( .A(n3082), .B(n4312), .Y(n1906) );
  NOR2BX1 U3740 ( .AN(n2285), .B(n352), .Y(n4312) );
  XNOR2X1 U3741 ( .A(n1280), .B(n1343), .Y(n2285) );
  CLKINVX1 U3742 ( .A(n3958), .Y(n3082) );
  XOR2X1 U3743 ( .A(n1407), .B(n1471), .Y(n3958) );
  XNOR2X1 U3744 ( .A(n3537), .B(n4313), .Y(n1891) );
  NOR2X1 U3745 ( .A(n2236), .B(n366), .Y(n4313) );
  XOR2X1 U3746 ( .A(n1290), .B(n1353), .Y(n2236) );
  CLKINVX1 U3747 ( .A(n3885), .Y(n3537) );
  XOR2X1 U3748 ( .A(n1417), .B(n1481), .Y(n3885) );
  XNOR2X1 U3749 ( .A(n3404), .B(n4314), .Y(n4223) );
  NOR2X1 U3750 ( .A(n346), .B(n3409), .Y(n4314) );
  XOR2X1 U3751 ( .A(n1297), .B(n1360), .Y(n3409) );
  XNOR2X1 U3752 ( .A(n1424), .B(n1488), .Y(n3404) );
  OAI222X1 U3753 ( .A0(n879), .A1(n4315), .B0(n905), .B1(n4316), .C0(n1203), 
        .C1(n854), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[101]) );
  XOR2X1 U3754 ( .A(n4228), .B(n4317), .Y(n4316) );
  XOR2X1 U3755 ( .A(n1897), .B(n1911), .Y(n4317) );
  XNOR2X1 U3756 ( .A(n3098), .B(n4318), .Y(n1911) );
  NOR2BX1 U3757 ( .AN(n2359), .B(n353), .Y(n4318) );
  XNOR2X1 U3758 ( .A(n1279), .B(n1342), .Y(n2359) );
  CLKINVX1 U3759 ( .A(n3968), .Y(n3098) );
  XOR2X1 U3760 ( .A(n1406), .B(n1470), .Y(n3968) );
  XNOR2X1 U3761 ( .A(n3556), .B(n4319), .Y(n1897) );
  NOR2X1 U3762 ( .A(n2242), .B(n367), .Y(n4319) );
  XOR2X1 U3763 ( .A(n1289), .B(n1352), .Y(n2242) );
  CLKINVX1 U3764 ( .A(n3895), .Y(n3556) );
  XOR2X1 U3765 ( .A(n1416), .B(n1480), .Y(n3895) );
  XNOR2X1 U3766 ( .A(n3424), .B(n4320), .Y(n4228) );
  NOR2BX1 U3767 ( .AN(n1551), .B(n3429), .Y(n4320) );
  XOR2X1 U3768 ( .A(n1296), .B(n1359), .Y(n3429) );
  XNOR2X1 U3769 ( .A(n1423), .B(n1487), .Y(n3424) );
  OAI222X1 U3770 ( .A0(n879), .A1(n4321), .B0(n904), .B1(n4322), .C0(n1204), 
        .C1(n856), .Y(Inst_AEAD_u_cc_u_cc_dp_istate[100]) );
  XOR2X1 U3771 ( .A(n4235), .B(n4323), .Y(n4322) );
  XOR2X1 U3772 ( .A(n1903), .B(n1916), .Y(n4323) );
  XNOR2X1 U3773 ( .A(n3109), .B(n4324), .Y(n1916) );
  NOR2X1 U3774 ( .A(n2425), .B(n368), .Y(n4324) );
  XOR2X1 U3775 ( .A(n1278), .B(n1341), .Y(n2425) );
  CLKINVX1 U3776 ( .A(n3975), .Y(n3109) );
  XOR2X1 U3777 ( .A(n1405), .B(n1469), .Y(n3975) );
  XNOR2X1 U3778 ( .A(n3576), .B(n4325), .Y(n1903) );
  NOR2X1 U3779 ( .A(n2251), .B(n369), .Y(n4325) );
  XOR2X1 U3780 ( .A(n1288), .B(n1351), .Y(n2251) );
  CLKINVX1 U3781 ( .A(n3902), .Y(n3576) );
  XOR2X1 U3782 ( .A(n1415), .B(n1479), .Y(n3902) );
  XNOR2X1 U3783 ( .A(n3444), .B(n4326), .Y(n4235) );
  NOR2X1 U3784 ( .A(n347), .B(n3449), .Y(n4326) );
  XOR2X1 U3785 ( .A(n1295), .B(n1358), .Y(n3449) );
  XNOR2X1 U3786 ( .A(n1422), .B(n1486), .Y(n3444) );
  OAI222X1 U3787 ( .A0(n879), .A1(n4327), .B0(n4328), .B1(n907), .C0(
        Inst_AEAD_u_input_n321), .C1(n855), .Y(
        Inst_AEAD_u_cc_u_cc_dp_istate[0]) );
  XOR2X1 U3788 ( .A(n4329), .B(n2233), .Y(n4328) );
  MXI2X1 U3789 ( .A(n2704), .B(n3675), .S0(n1474), .Y(n2233) );
  XOR2X1 U3790 ( .A(n1283), .B(n1346), .Y(n3675) );
  XOR2X1 U3791 ( .A(n1346), .B(n370), .Y(n2704) );
  XOR2X1 U3792 ( .A(n1979), .B(n2151), .Y(n4329) );
  MXI2X1 U3793 ( .A(n2902), .B(n4330), .S0(n1433), .Y(n2151) );
  CLKINVX1 U3794 ( .A(n2905), .Y(n4330) );
  XOR2X1 U3795 ( .A(n1241), .B(n378), .Y(n2905) );
  XNOR2X1 U3796 ( .A(n1241), .B(n1497), .Y(n2902) );
  MXI2X1 U3797 ( .A(n4232), .B(n2779), .S0(n341), .Y(n1979) );
  CLKINVX1 U3798 ( .A(n2784), .Y(n2779) );
  XNOR2X1 U3799 ( .A(n1312), .B(n350), .Y(n2784) );
  CLKINVX1 U3800 ( .A(n2783), .Y(n4232) );
  XOR2X1 U3801 ( .A(n1249), .B(n441), .Y(n2783) );
  MXI2X1 U3802 ( .A(n4331), .B(n4332), .S0(Inst_AEAD_u_cc_u_cc_ctrl_n37), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n123) );
  NAND3XL U3803 ( .A(n4333), .B(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), .C(
        Inst_AEAD_u_cc_u_cc_ctrl_round_2_), .Y(n4332) );
  AOI21X1 U3804 ( .A0(n4334), .A1(n4335), .B0(n4336), .Y(n4331) );
  MXI2X1 U3805 ( .A(n4337), .B(n4338), .S0(Inst_AEAD_u_cc_sel_tag[0]), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n122) );
  CLKNAND2X2 U3806 ( .A(n4334), .B(n4338), .Y(n4337) );
  MXI2X1 U3807 ( .A(n4339), .B(n4340), .S0(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), 
        .Y(Inst_AEAD_u_cc_u_cc_ctrl_n121) );
  MXI2X1 U3808 ( .A(n4341), .B(n4342), .S0(n4335), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n120) );
  CLKNAND2X2 U3809 ( .A(n4333), .B(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), .Y(
        n4342) );
  CLKINVX1 U3810 ( .A(n4339), .Y(n4333) );
  NAND3XL U3811 ( .A(Inst_AEAD_u_cc_sel_tag[0]), .B(n4338), .C(n4334), .Y(
        n4339) );
  CLKINVX1 U3812 ( .A(n4336), .Y(n4341) );
  OAI21X1 U3813 ( .A0(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), .A1(n4343), .B0(
        n4340), .Y(n4336) );
  OA21X1 U3814 ( .A0(Inst_AEAD_u_cc_sel_tag[0]), .A1(n4343), .B0(n4338), .Y(
        n4340) );
  CLKNAND2X2 U3815 ( .A(n4334), .B(n1626), .Y(n4338) );
  NOR4BX1 U3816 ( .AN(n4344), .B(n4345), .C(n997), .D(Inst_AEAD_u_cc_en_cmp), 
        .Y(n1626) );
  CLKINVX1 U3817 ( .A(n4334), .Y(n4343) );
  NOR2X1 U3818 ( .A(n1627), .B(rst), .Y(n4334) );
  CLKINVX1 U3819 ( .A(n1840), .Y(n1627) );
  AOI211X1 U3820 ( .A0(n4346), .A1(n997), .B0(n1609), .C0(n4347), .Y(n1840) );
  NOR2BX1 U3821 ( .AN(n4348), .B(n1605), .Y(n5081) );
  CLKINVX1 U3822 ( .A(n4349), .Y(n4346) );
  NOR2X1 U3823 ( .A(n4350), .B(n4351), .Y(Inst_AEAD_u_cc_u_cc_ctrl_n119) );
  AOI2BB1X1 U3824 ( .A0N(n4352), .A1N(n4353), .B0(n905), .Y(n4350) );
  CLKNAND2X2 U3825 ( .A(n853), .B(n873), .Y(n1857) );
  OAI22X1 U3826 ( .A0(n4354), .A1(n4355), .B0(n4356), .B1(n4351), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n118) );
  CLKINVX1 U3827 ( .A(n4357), .Y(n4351) );
  AOI221XL U3828 ( .A0(Inst_AEAD_u_cc_u_cc_ctrl_state_0_), .A1(n4358), .B0(
        n1609), .B1(Inst_AEAD_key_update), .C0(n4359), .Y(n4356) );
  OAI31X1 U3829 ( .A0(n4360), .A1(n4361), .A2(n4362), .B0(n338), .Y(n4359) );
  XNOR2X1 U3830 ( .A(n4335), .B(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_2_), .Y(n4362)
         );
  XOR2X1 U3831 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_1_), .Y(n4361) );
  NAND3XL U3832 ( .A(Inst_AEAD_u_cc_sel_tag[0]), .B(n4363), .C(n4345), .Y(
        n4360) );
  XOR2X1 U3833 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_3_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_n37), .Y(n4363) );
  OAI2B1X1 U3834 ( .A1N(n4347), .A0(n4364), .B0(n4353), .Y(n4358) );
  AOI211X1 U3835 ( .A0(n4349), .A1(n4365), .B0(n4366), .C0(n4345), .Y(n4353)
         );
  OAI21X1 U3836 ( .A0(n4354), .A1(n4367), .B0(n4368), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n117) );
  OAI31X1 U3837 ( .A0(n4369), .A1(n4370), .A2(n4366), .B0(n4357), .Y(n4368) );
  AOI211X1 U3838 ( .A0(n4371), .A1(n5073), .B0(rst), .C0(n4372), .Y(n4357) );
  AOI211X1 U3839 ( .A0(Inst_AEAD_bdo_ready), .A1(Inst_AEAD_u_cc_u_cc_ctrl_n52), 
        .B0(n4373), .C0(n1773), .Y(n4366) );
  OAI21X1 U3840 ( .A0(n1605), .A1(n4349), .B0(n4374), .Y(n4369) );
  NAND4X1 U3841 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_round_1_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_n37), .C(Inst_AEAD_u_cc_sel_tag[0]), .D(n4335), .Y(n4349) );
  CLKINVX1 U3842 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_round_2_), .Y(n4335) );
  AOI22XL U3843 ( .A0(n981), .A1(n4372), .B0(n4371), .B1(n5073), .Y(n4354) );
  OAI22X1 U3844 ( .A0(n4348), .A1(n1605), .B0(Inst_AEAD_bdi_valid), .B1(n4374), 
        .Y(n4372) );
  AOI2BB1X1 U3845 ( .A0N(Inst_AEAD_key_update), .A1N(n4375), .B0(n470), .Y(
        n4374) );
  NOR3X1 U3846 ( .A(n1639), .B(Inst_AEAD_u_input_ss_0_), .C(n1604), .Y(n4348)
         );
  CLKINVX1 U3847 ( .A(sdi_valid), .Y(n1604) );
  CLKINVX1 U3848 ( .A(Inst_AEAD_u_input_ss_1_), .Y(n1639) );
  MX2X1 U3849 ( .A(n856), .B(Inst_AEAD_u_cc_u_cc_ctrl_is_init_dat), .S0(n4376), 
        .Y(Inst_AEAD_u_cc_u_cc_ctrl_n116) );
  AOI21X1 U3850 ( .A0(n4377), .A1(n981), .B0(n5073), .Y(n4376) );
  NOR2X1 U3851 ( .A(n853), .B(rst), .Y(n5073) );
  OAI2B1X1 U3852 ( .A1N(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_1_), .A0(n4378), .B0(
        n4379), .Y(Inst_AEAD_u_cc_u_cc_ctrl_n115) );
  AO21X1 U3853 ( .A0(n4379), .A1(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_2_), .B0(
        n4378), .Y(Inst_AEAD_u_cc_u_cc_ctrl_n114) );
  OAI2B1X1 U3854 ( .A1N(Inst_AEAD_u_cc_u_cc_ctrl_rndcmp_3_), .A0(n4378), .B0(
        n4379), .Y(Inst_AEAD_u_cc_u_cc_ctrl_n113) );
  CLKNAND2X2 U3855 ( .A(n981), .B(n1839), .Y(n4379) );
  NAND3XL U3856 ( .A(n1605), .B(n937), .C(n4375), .Y(n1839) );
  CLKINVX1 U3857 ( .A(n4365), .Y(n1605) );
  NOR3X1 U3858 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .C(n4355), .Y(n4365) );
  CLKINVX1 U3859 ( .A(rst), .Y(n5077) );
  AOI211X1 U3860 ( .A0(n4380), .A1(Inst_AEAD_bdi_eot), .B0(rst), .C0(n4381), 
        .Y(n4378) );
  AOI31X1 U3861 ( .A0(n4375), .A1(n937), .A2(n4382), .B0(rst), .Y(
        Inst_AEAD_u_cc_u_cc_ctrl_n112) );
  CLKNAND2X2 U3862 ( .A(Inst_AEAD_u_cc_sel_key_lo), .B(n4381), .Y(n4382) );
  CLKINVX1 U3863 ( .A(Inst_AEAD_bdi_eot), .Y(n1763) );
  CLKINVX1 U3864 ( .A(n1609), .Y(n4375) );
  NOR3X1 U3865 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .C(
        Inst_AEAD_u_cc_u_cc_ctrl_state_0_), .Y(n1609) );
  OR3X1 U3866 ( .A(n868), .B(n1776), .C(n4345), .Y(Inst_AEAD_u_cc_en_state) );
  NOR3X1 U3867 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_0_), .B(
        Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .C(n4352), .Y(n4345) );
  NOR3X1 U3868 ( .A(n4355), .B(Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .C(n4367), 
        .Y(n1775) );
  CLKINVX1 U3869 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .Y(n4367) );
  AND2X1 U3870 ( .A(n4370), .B(n4373), .Y(Inst_AEAD_u_cc_en_cmp) );
  NOR2BX1 U3871 ( .AN(Inst_AEAD_u_cc_u_cc_dp_N712), .B(n1561), .Y(
        Inst_AEAD_msg_auth_valid) );
  NOR4X1 U3872 ( .A(n4383), .B(n4384), .C(n4385), .D(n4386), .Y(
        Inst_AEAD_u_cc_u_cc_dp_N712) );
  NAND4X1 U3873 ( .A(n4387), .B(n4388), .C(n4389), .D(n4390), .Y(n4386) );
  NOR4X1 U3874 ( .A(n4391), .B(n4392), .C(n4393), .D(n4394), .Y(n4390) );
  XNOR2X1 U3875 ( .A(Inst_AEAD_u_input_n320), .B(Inst_AEAD_bdo[1]), .Y(n4394)
         );
  XNOR2X1 U3876 ( .A(Inst_AEAD_u_input_n308), .B(Inst_AEAD_bdo[14]), .Y(n4393)
         );
  XNOR2X1 U3877 ( .A(Inst_AEAD_u_input_n309), .B(Inst_AEAD_bdo[13]), .Y(n4392)
         );
  XNOR2X1 U3878 ( .A(Inst_AEAD_u_input_n310), .B(Inst_AEAD_bdo[12]), .Y(n4391)
         );
  NOR4X1 U3879 ( .A(n4395), .B(n4396), .C(n4397), .D(n4398), .Y(n4389) );
  XNOR2X1 U3880 ( .A(Inst_AEAD_u_input_n316), .B(Inst_AEAD_bdo[5]), .Y(n4398)
         );
  XNOR2X1 U3881 ( .A(Inst_AEAD_u_input_n317), .B(Inst_AEAD_bdo[4]), .Y(n4397)
         );
  XNOR2X1 U3882 ( .A(Inst_AEAD_u_input_n318), .B(Inst_AEAD_bdo[3]), .Y(n4396)
         );
  XNOR2X1 U3883 ( .A(Inst_AEAD_u_input_n319), .B(Inst_AEAD_bdo[2]), .Y(n4395)
         );
  NOR4X1 U3884 ( .A(n4399), .B(n4400), .C(n4401), .D(n4402), .Y(n4388) );
  XNOR2X1 U3885 ( .A(Inst_AEAD_u_input_n313), .B(Inst_AEAD_bdo[9]), .Y(n4402)
         );
  XNOR2X1 U3886 ( .A(Inst_AEAD_u_input_n314), .B(Inst_AEAD_bdo[8]), .Y(n4401)
         );
  XNOR2X1 U3887 ( .A(Inst_AEAD_u_input_n315), .B(Inst_AEAD_bdo[6]), .Y(n4400)
         );
  XNOR2X1 U3888 ( .A(n1600), .B(Inst_AEAD_bdo[63]), .Y(n4399) );
  NOR4X1 U3889 ( .A(n4403), .B(n4404), .C(n4405), .D(n4406), .Y(n4387) );
  XNOR2X1 U3890 ( .A(Inst_AEAD_u_input_n304), .B(Inst_AEAD_bdo[30]), .Y(n4406)
         );
  XNOR2X1 U3891 ( .A(Inst_AEAD_u_input_n305), .B(Inst_AEAD_bdo[29]), .Y(n4405)
         );
  XNOR2X1 U3892 ( .A(Inst_AEAD_u_input_n306), .B(Inst_AEAD_bdo[28]), .Y(n4404)
         );
  XNOR2X1 U3893 ( .A(Inst_AEAD_u_input_n307), .B(Inst_AEAD_bdo[25]), .Y(n4403)
         );
  NAND4X1 U3894 ( .A(n4407), .B(n4408), .C(n4409), .D(n4410), .Y(n4385) );
  NOR4X1 U3895 ( .A(n4411), .B(n4412), .C(n4413), .D(n4414), .Y(n4410) );
  XNOR2X1 U3896 ( .A(Inst_AEAD_bdo[17]), .B(n1716), .Y(n4414) );
  XNOR2X1 U3897 ( .A(Inst_AEAD_bdo[16]), .B(n1715), .Y(n4413) );
  XNOR2X1 U3898 ( .A(Inst_AEAD_bdo[15]), .B(n2669), .Y(n4412) );
  XNOR2X1 U3899 ( .A(Inst_AEAD_bdo[7]), .B(n1976), .Y(n4411) );
  NOR4X1 U3900 ( .A(n4415), .B(n4416), .C(n4417), .D(n4418), .Y(n4409) );
  XNOR2X1 U3901 ( .A(Inst_AEAD_bdo[21]), .B(n1720), .Y(n4418) );
  XNOR2X1 U3902 ( .A(Inst_AEAD_bdo[20]), .B(n1719), .Y(n4417) );
  XNOR2X1 U3903 ( .A(Inst_AEAD_bdo[19]), .B(n1718), .Y(n4416) );
  XNOR2X1 U3904 ( .A(Inst_AEAD_bdo[18]), .B(n1717), .Y(n4415) );
  NOR4X1 U3905 ( .A(n4419), .B(n4420), .C(n4421), .D(n4422), .Y(n4408) );
  XNOR2X1 U3906 ( .A(Inst_AEAD_bdo[26]), .B(n1725), .Y(n4422) );
  XNOR2X1 U3907 ( .A(Inst_AEAD_bdo[24]), .B(n1722), .Y(n4421) );
  XNOR2X1 U3908 ( .A(Inst_AEAD_bdo[23]), .B(n2595), .Y(n4420) );
  XNOR2X1 U3909 ( .A(Inst_AEAD_bdo[22]), .B(n1721), .Y(n4419) );
  NOR4X1 U3910 ( .A(n4423), .B(n4424), .C(n4425), .D(n4426), .Y(n4407) );
  XNOR2X1 U3911 ( .A(Inst_AEAD_u_input_n311), .B(Inst_AEAD_bdo[11]), .Y(n4426)
         );
  XNOR2X1 U3912 ( .A(Inst_AEAD_u_input_n312), .B(Inst_AEAD_bdo[10]), .Y(n4425)
         );
  XNOR2X1 U3913 ( .A(Inst_AEAD_u_input_n321), .B(Inst_AEAD_bdo[0]), .Y(n4424)
         );
  XNOR2X1 U3914 ( .A(Inst_AEAD_bdo[27]), .B(n1726), .Y(n4423) );
  NAND4X1 U3915 ( .A(n4427), .B(n4428), .C(n4429), .D(n4430), .Y(n4384) );
  NOR4X1 U3916 ( .A(n4431), .B(n4432), .C(n4433), .D(n4434), .Y(n4430) );
  XNOR2X1 U3917 ( .A(n1579), .B(Inst_AEAD_bdo[50]), .Y(n4434) );
  XNOR2X1 U3918 ( .A(n1580), .B(Inst_AEAD_bdo[49]), .Y(n4433) );
  XNOR2X1 U3919 ( .A(n1581), .B(Inst_AEAD_bdo[48]), .Y(n4432) );
  XNOR2X1 U3920 ( .A(n1602), .B(Inst_AEAD_bdo[47]), .Y(n4431) );
  NOR4X1 U3921 ( .A(n4435), .B(n4436), .C(n4437), .D(n4438), .Y(n4429) );
  XNOR2X1 U3922 ( .A(n1575), .B(Inst_AEAD_bdo[54]), .Y(n4438) );
  XNOR2X1 U3923 ( .A(n1576), .B(Inst_AEAD_bdo[53]), .Y(n4437) );
  XNOR2X1 U3924 ( .A(n1577), .B(Inst_AEAD_bdo[52]), .Y(n4436) );
  XNOR2X1 U3925 ( .A(n1578), .B(Inst_AEAD_bdo[51]), .Y(n4435) );
  NOR4X1 U3926 ( .A(n4439), .B(n4440), .C(n4441), .D(n4442), .Y(n4428) );
  XNOR2X1 U3927 ( .A(n1572), .B(Inst_AEAD_bdo[58]), .Y(n4442) );
  XNOR2X1 U3928 ( .A(n1573), .B(Inst_AEAD_bdo[57]), .Y(n4441) );
  XNOR2X1 U3929 ( .A(n1574), .B(Inst_AEAD_bdo[56]), .Y(n4440) );
  XNOR2X1 U3930 ( .A(n1601), .B(Inst_AEAD_bdo[55]), .Y(n4439) );
  NOR4X1 U3931 ( .A(n4443), .B(n4444), .C(n4445), .D(n4446), .Y(n4427) );
  XNOR2X1 U3932 ( .A(n1568), .B(Inst_AEAD_bdo[62]), .Y(n4446) );
  XNOR2X1 U3933 ( .A(n1569), .B(Inst_AEAD_bdo[61]), .Y(n4445) );
  XNOR2X1 U3934 ( .A(n1570), .B(Inst_AEAD_bdo[60]), .Y(n4444) );
  XNOR2X1 U3935 ( .A(n1571), .B(Inst_AEAD_bdo[59]), .Y(n4443) );
  NAND4X1 U3936 ( .A(n4447), .B(n4448), .C(n4449), .D(n4450), .Y(n4383) );
  NOR4X1 U3937 ( .A(n4451), .B(n4452), .C(n4453), .D(n4454), .Y(n4450) );
  XNOR2X1 U3938 ( .A(n1593), .B(Inst_AEAD_bdo[34]), .Y(n4454) );
  XNOR2X1 U3939 ( .A(n1594), .B(Inst_AEAD_bdo[33]), .Y(n4453) );
  XNOR2X1 U3940 ( .A(n1595), .B(Inst_AEAD_bdo[32]), .Y(n4452) );
  XNOR2X1 U3941 ( .A(Inst_AEAD_u_input_n303), .B(Inst_AEAD_bdo[31]), .Y(n4451)
         );
  NOR4X1 U3942 ( .A(n4455), .B(n4456), .C(n4457), .D(n4458), .Y(n4449) );
  XNOR2X1 U3943 ( .A(n1589), .B(Inst_AEAD_bdo[38]), .Y(n4458) );
  XNOR2X1 U3944 ( .A(n1590), .B(Inst_AEAD_bdo[37]), .Y(n4457) );
  XNOR2X1 U3945 ( .A(n1591), .B(Inst_AEAD_bdo[36]), .Y(n4456) );
  XNOR2X1 U3946 ( .A(n1592), .B(Inst_AEAD_bdo[35]), .Y(n4455) );
  NOR4X1 U3947 ( .A(n4459), .B(n4460), .C(n4461), .D(n4462), .Y(n4448) );
  XNOR2X1 U3948 ( .A(n1586), .B(Inst_AEAD_bdo[42]), .Y(n4462) );
  XNOR2X1 U3949 ( .A(n1587), .B(Inst_AEAD_bdo[41]), .Y(n4461) );
  XNOR2X1 U3950 ( .A(n1588), .B(Inst_AEAD_bdo[40]), .Y(n4460) );
  XNOR2X1 U3951 ( .A(n1603), .B(Inst_AEAD_bdo[39]), .Y(n4459) );
  NOR4X1 U3952 ( .A(n4463), .B(n4464), .C(n4465), .D(n4466), .Y(n4447) );
  XNOR2X1 U3953 ( .A(n1582), .B(Inst_AEAD_bdo[46]), .Y(n4466) );
  XNOR2X1 U3954 ( .A(n1583), .B(Inst_AEAD_bdo[45]), .Y(n4465) );
  XNOR2X1 U3955 ( .A(n1584), .B(Inst_AEAD_bdo[44]), .Y(n4464) );
  XNOR2X1 U3956 ( .A(n1585), .B(Inst_AEAD_bdo[43]), .Y(n4463) );
  NOR2BX1 U3957 ( .AN(n4373), .B(n1773), .Y(Inst_AEAD_msg_auth_done) );
  NOR2X1 U3958 ( .A(n4371), .B(Inst_AEAD_u_cc_u_cc_ctrl_n52), .Y(n4373) );
  NAND4X1 U3959 ( .A(n4467), .B(n4468), .C(n4469), .D(n4470), .Y(
        Inst_AEAD_key[9]) );
  MXI2X1 U3960 ( .A(n4471), .B(n4472), .S0(randd[41]), .Y(n4470) );
  OAI21X1 U3961 ( .A0(IDtReg[41]), .A1(n4473), .B0(n4474), .Y(n4472) );
  NOR2X1 U3962 ( .A(n4475), .B(n4473), .Y(n4471) );
  MXI2X1 U3963 ( .A(n4476), .B(n4477), .S0(randd[9]), .Y(n4469) );
  OAI21X1 U3964 ( .A0(IDtReg[9]), .A1(n4478), .B0(n4479), .Y(n4477) );
  NOR2X1 U3965 ( .A(n4480), .B(n4478), .Y(n4476) );
  MXI2X1 U3966 ( .A(n4481), .B(n4482), .S0(rand_in[41]), .Y(n4468) );
  OAI22X1 U3967 ( .A0(IDtReg[41]), .A1(n4483), .B0(IDstReg[41]), .B1(n4484), 
        .Y(n4482) );
  OAI2B2X1 U3968 ( .A1N(IDstReg[41]), .A0(n4484), .B0(n4475), .B1(n4483), .Y(
        n4481) );
  CLKINVX1 U3969 ( .A(IDtReg[41]), .Y(n4475) );
  MXI2X1 U3970 ( .A(n4485), .B(n4486), .S0(rand_in[9]), .Y(n4467) );
  OAI22X1 U3971 ( .A0(IDtReg[9]), .A1(n4487), .B0(IDstReg[9]), .B1(n4488), .Y(
        n4486) );
  OAI2B2X1 U3972 ( .A1N(IDstReg[9]), .A0(n4488), .B0(n4480), .B1(n4487), .Y(
        n4485) );
  CLKINVX1 U3973 ( .A(IDtReg[9]), .Y(n4480) );
  NAND4X1 U3974 ( .A(n4489), .B(n4490), .C(n4491), .D(n4492), .Y(
        Inst_AEAD_key[8]) );
  MXI2X1 U3975 ( .A(n4493), .B(n4494), .S0(randd[40]), .Y(n4492) );
  OAI21X1 U3976 ( .A0(IDtReg[40]), .A1(n4473), .B0(n4474), .Y(n4494) );
  NOR2X1 U3977 ( .A(n4495), .B(n4473), .Y(n4493) );
  MXI2X1 U3978 ( .A(n4496), .B(n4497), .S0(randd[8]), .Y(n4491) );
  OAI21X1 U3979 ( .A0(IDtReg[8]), .A1(n4478), .B0(n4479), .Y(n4497) );
  NOR2X1 U3980 ( .A(n4498), .B(n4478), .Y(n4496) );
  MXI2X1 U3981 ( .A(n4499), .B(n4500), .S0(rand_in[40]), .Y(n4490) );
  OAI22X1 U3982 ( .A0(IDtReg[40]), .A1(n4483), .B0(IDstReg[40]), .B1(n4484), 
        .Y(n4500) );
  OAI2B2X1 U3983 ( .A1N(IDstReg[40]), .A0(n4484), .B0(n4495), .B1(n4483), .Y(
        n4499) );
  CLKINVX1 U3984 ( .A(IDtReg[40]), .Y(n4495) );
  MXI2X1 U3985 ( .A(n4501), .B(n4502), .S0(rand_in[8]), .Y(n4489) );
  OAI22X1 U3986 ( .A0(IDtReg[8]), .A1(n4487), .B0(IDstReg[8]), .B1(n4488), .Y(
        n4502) );
  OAI2B2X1 U3987 ( .A1N(IDstReg[8]), .A0(n4488), .B0(n4498), .B1(n4487), .Y(
        n4501) );
  CLKINVX1 U3988 ( .A(IDtReg[8]), .Y(n4498) );
  NAND4X1 U3989 ( .A(n4503), .B(n4504), .C(n4505), .D(n4506), .Y(
        Inst_AEAD_key[7]) );
  MXI2X1 U3990 ( .A(n4507), .B(n4508), .S0(randd[39]), .Y(n4506) );
  OAI21X1 U3991 ( .A0(IDtReg[39]), .A1(n4473), .B0(n4474), .Y(n4508) );
  NOR2X1 U3992 ( .A(n4509), .B(n4473), .Y(n4507) );
  MXI2X1 U3993 ( .A(n4510), .B(n4511), .S0(randd[7]), .Y(n4505) );
  OAI21X1 U3994 ( .A0(IDtReg[7]), .A1(n4478), .B0(n4479), .Y(n4511) );
  NOR2X1 U3995 ( .A(n4512), .B(n4478), .Y(n4510) );
  MXI2X1 U3996 ( .A(n4513), .B(n4514), .S0(rand_in[39]), .Y(n4504) );
  OAI22X1 U3997 ( .A0(IDtReg[39]), .A1(n4483), .B0(IDstReg[39]), .B1(n4484), 
        .Y(n4514) );
  OAI2B2X1 U3998 ( .A1N(IDstReg[39]), .A0(n4484), .B0(n4509), .B1(n4483), .Y(
        n4513) );
  CLKINVX1 U3999 ( .A(IDtReg[39]), .Y(n4509) );
  MXI2X1 U4000 ( .A(n4515), .B(n4516), .S0(rand_in[7]), .Y(n4503) );
  OAI22X1 U4001 ( .A0(IDtReg[7]), .A1(n4487), .B0(IDstReg[7]), .B1(n4488), .Y(
        n4516) );
  OAI2B2X1 U4002 ( .A1N(IDstReg[7]), .A0(n4488), .B0(n4512), .B1(n4487), .Y(
        n4515) );
  CLKINVX1 U4003 ( .A(IDtReg[7]), .Y(n4512) );
  NAND4X1 U4004 ( .A(n4517), .B(n4518), .C(n4519), .D(n4520), .Y(
        Inst_AEAD_key[6]) );
  MXI2X1 U4005 ( .A(n4521), .B(n4522), .S0(randd[38]), .Y(n4520) );
  OAI21X1 U4006 ( .A0(IDtReg[38]), .A1(n4473), .B0(n4474), .Y(n4522) );
  NOR2X1 U4007 ( .A(n4523), .B(n4473), .Y(n4521) );
  MXI2X1 U4008 ( .A(n4524), .B(n4525), .S0(randd[6]), .Y(n4519) );
  OAI21X1 U4009 ( .A0(IDtReg[6]), .A1(n4478), .B0(n4479), .Y(n4525) );
  NOR2X1 U4010 ( .A(n4526), .B(n4478), .Y(n4524) );
  MXI2X1 U4011 ( .A(n4527), .B(n4528), .S0(rand_in[38]), .Y(n4518) );
  OAI22X1 U4012 ( .A0(IDtReg[38]), .A1(n4483), .B0(IDstReg[38]), .B1(n4484), 
        .Y(n4528) );
  OAI2B2X1 U4013 ( .A1N(IDstReg[38]), .A0(n4484), .B0(n4523), .B1(n4483), .Y(
        n4527) );
  CLKINVX1 U4014 ( .A(IDtReg[38]), .Y(n4523) );
  MXI2X1 U4015 ( .A(n4529), .B(n4530), .S0(rand_in[6]), .Y(n4517) );
  OAI22X1 U4016 ( .A0(IDtReg[6]), .A1(n4487), .B0(IDstReg[6]), .B1(n4488), .Y(
        n4530) );
  OAI2B2X1 U4017 ( .A1N(IDstReg[6]), .A0(n4488), .B0(n4526), .B1(n4487), .Y(
        n4529) );
  CLKINVX1 U4018 ( .A(IDtReg[6]), .Y(n4526) );
  NAND4X1 U4019 ( .A(n4531), .B(n4532), .C(n4533), .D(n4534), .Y(
        Inst_AEAD_key[5]) );
  MXI2X1 U4020 ( .A(n4535), .B(n4536), .S0(randd[37]), .Y(n4534) );
  OAI21X1 U4021 ( .A0(IDtReg[37]), .A1(n4473), .B0(n4474), .Y(n4536) );
  NOR2X1 U4022 ( .A(n4537), .B(n4473), .Y(n4535) );
  MXI2X1 U4023 ( .A(n4538), .B(n4539), .S0(randd[5]), .Y(n4533) );
  OAI21X1 U4024 ( .A0(IDtReg[5]), .A1(n4478), .B0(n4479), .Y(n4539) );
  NOR2X1 U4025 ( .A(n4540), .B(n4478), .Y(n4538) );
  MXI2X1 U4026 ( .A(n4541), .B(n4542), .S0(rand_in[37]), .Y(n4532) );
  OAI22X1 U4027 ( .A0(IDtReg[37]), .A1(n4483), .B0(IDstReg[37]), .B1(n4484), 
        .Y(n4542) );
  OAI2B2X1 U4028 ( .A1N(IDstReg[37]), .A0(n4484), .B0(n4537), .B1(n4483), .Y(
        n4541) );
  CLKINVX1 U4029 ( .A(IDtReg[37]), .Y(n4537) );
  MXI2X1 U4030 ( .A(n4543), .B(n4544), .S0(rand_in[5]), .Y(n4531) );
  OAI22X1 U4031 ( .A0(IDtReg[5]), .A1(n4487), .B0(IDstReg[5]), .B1(n4488), .Y(
        n4544) );
  OAI2B2X1 U4032 ( .A1N(IDstReg[5]), .A0(n4488), .B0(n4540), .B1(n4487), .Y(
        n4543) );
  CLKINVX1 U4033 ( .A(IDtReg[5]), .Y(n4540) );
  NAND4X1 U4034 ( .A(n4545), .B(n4546), .C(n4547), .D(n4548), .Y(
        Inst_AEAD_key[4]) );
  MXI2X1 U4035 ( .A(n4549), .B(n4550), .S0(randd[36]), .Y(n4548) );
  OAI21X1 U4036 ( .A0(IDtReg[36]), .A1(n4473), .B0(n4474), .Y(n4550) );
  NOR2X1 U4037 ( .A(n4551), .B(n4473), .Y(n4549) );
  MXI2X1 U4038 ( .A(n4552), .B(n4553), .S0(randd[4]), .Y(n4547) );
  OAI21X1 U4039 ( .A0(IDtReg[4]), .A1(n4478), .B0(n4479), .Y(n4553) );
  NOR2X1 U4040 ( .A(n4554), .B(n4478), .Y(n4552) );
  MXI2X1 U4041 ( .A(n4555), .B(n4556), .S0(rand_in[36]), .Y(n4546) );
  OAI22X1 U4042 ( .A0(IDtReg[36]), .A1(n4483), .B0(IDstReg[36]), .B1(n4484), 
        .Y(n4556) );
  OAI2B2X1 U4043 ( .A1N(IDstReg[36]), .A0(n4484), .B0(n4551), .B1(n4483), .Y(
        n4555) );
  CLKINVX1 U4044 ( .A(IDtReg[36]), .Y(n4551) );
  MXI2X1 U4045 ( .A(n4557), .B(n4558), .S0(rand_in[4]), .Y(n4545) );
  OAI22X1 U4046 ( .A0(IDtReg[4]), .A1(n4487), .B0(IDstReg[4]), .B1(n4488), .Y(
        n4558) );
  OAI2B2X1 U4047 ( .A1N(IDstReg[4]), .A0(n4488), .B0(n4554), .B1(n4487), .Y(
        n4557) );
  CLKINVX1 U4048 ( .A(IDtReg[4]), .Y(n4554) );
  NAND4X1 U4049 ( .A(n4559), .B(n4560), .C(n4561), .D(n4562), .Y(
        Inst_AEAD_key[3]) );
  MXI2X1 U4050 ( .A(n4563), .B(n4564), .S0(randd[35]), .Y(n4562) );
  OAI21X1 U4051 ( .A0(IDtReg[35]), .A1(n4473), .B0(n4474), .Y(n4564) );
  NOR2X1 U4052 ( .A(n4565), .B(n4473), .Y(n4563) );
  MXI2X1 U4053 ( .A(n4566), .B(n4567), .S0(randd[3]), .Y(n4561) );
  OAI21X1 U4054 ( .A0(IDtReg[3]), .A1(n4478), .B0(n4479), .Y(n4567) );
  NOR2X1 U4055 ( .A(n4568), .B(n4478), .Y(n4566) );
  MXI2X1 U4056 ( .A(n4569), .B(n4570), .S0(rand_in[35]), .Y(n4560) );
  OAI22X1 U4057 ( .A0(IDtReg[35]), .A1(n4483), .B0(IDstReg[35]), .B1(n4484), 
        .Y(n4570) );
  OAI2B2X1 U4058 ( .A1N(IDstReg[35]), .A0(n4484), .B0(n4565), .B1(n4483), .Y(
        n4569) );
  CLKINVX1 U4059 ( .A(IDtReg[35]), .Y(n4565) );
  MXI2X1 U4060 ( .A(n4571), .B(n4572), .S0(rand_in[3]), .Y(n4559) );
  OAI22X1 U4061 ( .A0(IDtReg[3]), .A1(n4487), .B0(IDstReg[3]), .B1(n4488), .Y(
        n4572) );
  OAI2B2X1 U4062 ( .A1N(IDstReg[3]), .A0(n4488), .B0(n4568), .B1(n4487), .Y(
        n4571) );
  CLKINVX1 U4063 ( .A(IDtReg[3]), .Y(n4568) );
  NAND4X1 U4064 ( .A(n4573), .B(n4574), .C(n4575), .D(n4576), .Y(
        Inst_AEAD_key[31]) );
  MXI2X1 U4065 ( .A(n4577), .B(n4578), .S0(randd[63]), .Y(n4576) );
  OAI21X1 U4066 ( .A0(IDtReg[63]), .A1(n4473), .B0(n4474), .Y(n4578) );
  NOR2X1 U4067 ( .A(n4579), .B(n4473), .Y(n4577) );
  MXI2X1 U4068 ( .A(n4580), .B(n4581), .S0(randd[31]), .Y(n4575) );
  OAI21X1 U4069 ( .A0(IDtReg[31]), .A1(n4478), .B0(n4479), .Y(n4581) );
  NOR2X1 U4070 ( .A(n4582), .B(n4478), .Y(n4580) );
  MXI2X1 U4071 ( .A(n4583), .B(n4584), .S0(rand_in[31]), .Y(n4574) );
  OAI22X1 U4072 ( .A0(IDtReg[31]), .A1(n4487), .B0(IDstReg[31]), .B1(n4488), 
        .Y(n4584) );
  OAI2B2X1 U4073 ( .A1N(IDstReg[31]), .A0(n4488), .B0(n4582), .B1(n4487), .Y(
        n4583) );
  CLKINVX1 U4074 ( .A(IDtReg[31]), .Y(n4582) );
  MXI2X1 U4075 ( .A(n4585), .B(n4586), .S0(rand_in[63]), .Y(n4573) );
  OAI22X1 U4076 ( .A0(IDtReg[63]), .A1(n4483), .B0(IDstReg[63]), .B1(n4484), 
        .Y(n4586) );
  OAI2B2X1 U4077 ( .A1N(IDstReg[63]), .A0(n4484), .B0(n4579), .B1(n4483), .Y(
        n4585) );
  CLKINVX1 U4078 ( .A(IDtReg[63]), .Y(n4579) );
  NAND4X1 U4079 ( .A(n4587), .B(n4588), .C(n4589), .D(n4590), .Y(
        Inst_AEAD_key[30]) );
  MXI2X1 U4080 ( .A(n4591), .B(n4592), .S0(randd[62]), .Y(n4590) );
  OAI21X1 U4081 ( .A0(IDtReg[62]), .A1(n4473), .B0(n4474), .Y(n4592) );
  NOR2X1 U4082 ( .A(n4593), .B(n4473), .Y(n4591) );
  MXI2X1 U4083 ( .A(n4594), .B(n4595), .S0(randd[30]), .Y(n4589) );
  OAI21X1 U4084 ( .A0(IDtReg[30]), .A1(n4478), .B0(n4479), .Y(n4595) );
  NOR2X1 U4085 ( .A(n4596), .B(n4478), .Y(n4594) );
  MXI2X1 U4086 ( .A(n4597), .B(n4598), .S0(rand_in[30]), .Y(n4588) );
  OAI22X1 U4087 ( .A0(IDtReg[30]), .A1(n4487), .B0(IDstReg[30]), .B1(n4488), 
        .Y(n4598) );
  OAI2B2X1 U4088 ( .A1N(IDstReg[30]), .A0(n4488), .B0(n4596), .B1(n4487), .Y(
        n4597) );
  CLKINVX1 U4089 ( .A(IDtReg[30]), .Y(n4596) );
  MXI2X1 U4090 ( .A(n4599), .B(n4600), .S0(rand_in[62]), .Y(n4587) );
  OAI22X1 U4091 ( .A0(IDtReg[62]), .A1(n4483), .B0(IDstReg[62]), .B1(n4484), 
        .Y(n4600) );
  OAI2B2X1 U4092 ( .A1N(IDstReg[62]), .A0(n4484), .B0(n4593), .B1(n4483), .Y(
        n4599) );
  CLKINVX1 U4093 ( .A(IDtReg[62]), .Y(n4593) );
  NAND4X1 U4094 ( .A(n4601), .B(n4602), .C(n4603), .D(n4604), .Y(
        Inst_AEAD_key[2]) );
  MXI2X1 U4095 ( .A(n4605), .B(n4606), .S0(randd[34]), .Y(n4604) );
  OAI21X1 U4096 ( .A0(IDtReg[34]), .A1(n4473), .B0(n4474), .Y(n4606) );
  NOR2X1 U4097 ( .A(n4607), .B(n4473), .Y(n4605) );
  MXI2X1 U4098 ( .A(n4608), .B(n4609), .S0(randd[2]), .Y(n4603) );
  OAI21X1 U4099 ( .A0(IDtReg[2]), .A1(n4478), .B0(n4479), .Y(n4609) );
  NOR2X1 U4100 ( .A(n4610), .B(n4478), .Y(n4608) );
  MXI2X1 U4101 ( .A(n4611), .B(n4612), .S0(rand_in[2]), .Y(n4602) );
  OAI22X1 U4102 ( .A0(IDtReg[2]), .A1(n4487), .B0(IDstReg[2]), .B1(n4488), .Y(
        n4612) );
  OAI2B2X1 U4103 ( .A1N(IDstReg[2]), .A0(n4488), .B0(n4610), .B1(n4487), .Y(
        n4611) );
  CLKINVX1 U4104 ( .A(IDtReg[2]), .Y(n4610) );
  MXI2X1 U4105 ( .A(n4613), .B(n4614), .S0(rand_in[34]), .Y(n4601) );
  OAI22X1 U4106 ( .A0(IDtReg[34]), .A1(n4483), .B0(IDstReg[34]), .B1(n4484), 
        .Y(n4614) );
  OAI2B2X1 U4107 ( .A1N(IDstReg[34]), .A0(n4484), .B0(n4607), .B1(n4483), .Y(
        n4613) );
  CLKINVX1 U4108 ( .A(IDtReg[34]), .Y(n4607) );
  NAND4X1 U4109 ( .A(n4615), .B(n4616), .C(n4617), .D(n4618), .Y(
        Inst_AEAD_key[29]) );
  MXI2X1 U4110 ( .A(n4619), .B(n4620), .S0(randd[61]), .Y(n4618) );
  OAI21X1 U4111 ( .A0(IDtReg[61]), .A1(n4473), .B0(n4474), .Y(n4620) );
  NOR2X1 U4112 ( .A(n4621), .B(n4473), .Y(n4619) );
  MXI2X1 U4113 ( .A(n4622), .B(n4623), .S0(randd[29]), .Y(n4617) );
  OAI21X1 U4114 ( .A0(IDtReg[29]), .A1(n4478), .B0(n4479), .Y(n4623) );
  NOR2X1 U4115 ( .A(n4624), .B(n4478), .Y(n4622) );
  MXI2X1 U4116 ( .A(n4625), .B(n4626), .S0(rand_in[29]), .Y(n4616) );
  OAI22X1 U4117 ( .A0(IDtReg[29]), .A1(n4487), .B0(IDstReg[29]), .B1(n4488), 
        .Y(n4626) );
  OAI2B2X1 U4118 ( .A1N(IDstReg[29]), .A0(n4488), .B0(n4624), .B1(n4487), .Y(
        n4625) );
  CLKINVX1 U4119 ( .A(IDtReg[29]), .Y(n4624) );
  MXI2X1 U4120 ( .A(n4627), .B(n4628), .S0(rand_in[61]), .Y(n4615) );
  OAI22X1 U4121 ( .A0(IDtReg[61]), .A1(n4483), .B0(IDstReg[61]), .B1(n4484), 
        .Y(n4628) );
  OAI2B2X1 U4122 ( .A1N(IDstReg[61]), .A0(n4484), .B0(n4621), .B1(n4483), .Y(
        n4627) );
  CLKINVX1 U4123 ( .A(IDtReg[61]), .Y(n4621) );
  NAND4X1 U4124 ( .A(n4629), .B(n4630), .C(n4631), .D(n4632), .Y(
        Inst_AEAD_key[28]) );
  MXI2X1 U4125 ( .A(n4633), .B(n4634), .S0(randd[60]), .Y(n4632) );
  OAI21X1 U4126 ( .A0(IDtReg[60]), .A1(n4473), .B0(n4474), .Y(n4634) );
  NOR2X1 U4127 ( .A(n4635), .B(n4473), .Y(n4633) );
  MXI2X1 U4128 ( .A(n4636), .B(n4637), .S0(randd[28]), .Y(n4631) );
  OAI21X1 U4129 ( .A0(IDtReg[28]), .A1(n4478), .B0(n4479), .Y(n4637) );
  NOR2X1 U4130 ( .A(n4638), .B(n4478), .Y(n4636) );
  MXI2X1 U4131 ( .A(n4639), .B(n4640), .S0(rand_in[28]), .Y(n4630) );
  OAI22X1 U4132 ( .A0(IDtReg[28]), .A1(n4487), .B0(IDstReg[28]), .B1(n4488), 
        .Y(n4640) );
  OAI2B2X1 U4133 ( .A1N(IDstReg[28]), .A0(n4488), .B0(n4638), .B1(n4487), .Y(
        n4639) );
  CLKINVX1 U4134 ( .A(IDtReg[28]), .Y(n4638) );
  MXI2X1 U4135 ( .A(n4641), .B(n4642), .S0(rand_in[60]), .Y(n4629) );
  OAI22X1 U4136 ( .A0(IDtReg[60]), .A1(n4483), .B0(IDstReg[60]), .B1(n4484), 
        .Y(n4642) );
  OAI2B2X1 U4137 ( .A1N(IDstReg[60]), .A0(n4484), .B0(n4635), .B1(n4483), .Y(
        n4641) );
  CLKINVX1 U4138 ( .A(IDtReg[60]), .Y(n4635) );
  NAND4X1 U4139 ( .A(n4643), .B(n4644), .C(n4645), .D(n4646), .Y(
        Inst_AEAD_key[27]) );
  MXI2X1 U4140 ( .A(n4647), .B(n4648), .S0(randd[59]), .Y(n4646) );
  OAI21X1 U4141 ( .A0(IDtReg[59]), .A1(n4473), .B0(n4474), .Y(n4648) );
  NOR2X1 U4142 ( .A(n4649), .B(n4473), .Y(n4647) );
  MXI2X1 U4143 ( .A(n4650), .B(n4651), .S0(randd[27]), .Y(n4645) );
  OAI21X1 U4144 ( .A0(IDtReg[27]), .A1(n4478), .B0(n4479), .Y(n4651) );
  NOR2X1 U4145 ( .A(n4652), .B(n4478), .Y(n4650) );
  MXI2X1 U4146 ( .A(n4653), .B(n4654), .S0(rand_in[27]), .Y(n4644) );
  OAI22X1 U4147 ( .A0(IDtReg[27]), .A1(n4487), .B0(IDstReg[27]), .B1(n4488), 
        .Y(n4654) );
  OAI2B2X1 U4148 ( .A1N(IDstReg[27]), .A0(n4488), .B0(n4652), .B1(n4487), .Y(
        n4653) );
  CLKINVX1 U4149 ( .A(IDtReg[27]), .Y(n4652) );
  MXI2X1 U4150 ( .A(n4655), .B(n4656), .S0(rand_in[59]), .Y(n4643) );
  OAI22X1 U4151 ( .A0(IDtReg[59]), .A1(n4483), .B0(IDstReg[59]), .B1(n4484), 
        .Y(n4656) );
  OAI2B2X1 U4152 ( .A1N(IDstReg[59]), .A0(n4484), .B0(n4649), .B1(n4483), .Y(
        n4655) );
  CLKINVX1 U4153 ( .A(IDtReg[59]), .Y(n4649) );
  NAND4X1 U4154 ( .A(n4657), .B(n4658), .C(n4659), .D(n4660), .Y(
        Inst_AEAD_key[26]) );
  MXI2X1 U4155 ( .A(n4661), .B(n4662), .S0(randd[58]), .Y(n4660) );
  OAI21X1 U4156 ( .A0(IDtReg[58]), .A1(n4473), .B0(n4474), .Y(n4662) );
  NOR2X1 U4157 ( .A(n4663), .B(n4473), .Y(n4661) );
  MXI2X1 U4158 ( .A(n4664), .B(n4665), .S0(randd[26]), .Y(n4659) );
  OAI21X1 U4159 ( .A0(IDtReg[26]), .A1(n4478), .B0(n4479), .Y(n4665) );
  NOR2X1 U4160 ( .A(n4666), .B(n4478), .Y(n4664) );
  MXI2X1 U4161 ( .A(n4667), .B(n4668), .S0(rand_in[26]), .Y(n4658) );
  OAI22X1 U4162 ( .A0(IDtReg[26]), .A1(n4487), .B0(IDstReg[26]), .B1(n4488), 
        .Y(n4668) );
  OAI2B2X1 U4163 ( .A1N(IDstReg[26]), .A0(n4488), .B0(n4666), .B1(n4487), .Y(
        n4667) );
  CLKINVX1 U4164 ( .A(IDtReg[26]), .Y(n4666) );
  MXI2X1 U4165 ( .A(n4669), .B(n4670), .S0(rand_in[58]), .Y(n4657) );
  OAI22X1 U4166 ( .A0(IDtReg[58]), .A1(n4483), .B0(IDstReg[58]), .B1(n4484), 
        .Y(n4670) );
  OAI2B2X1 U4167 ( .A1N(IDstReg[58]), .A0(n4484), .B0(n4663), .B1(n4483), .Y(
        n4669) );
  CLKINVX1 U4168 ( .A(IDtReg[58]), .Y(n4663) );
  NAND4X1 U4169 ( .A(n4671), .B(n4672), .C(n4673), .D(n4674), .Y(
        Inst_AEAD_key[25]) );
  MXI2X1 U4170 ( .A(n4675), .B(n4676), .S0(randd[57]), .Y(n4674) );
  OAI21X1 U4171 ( .A0(IDtReg[57]), .A1(n4473), .B0(n4474), .Y(n4676) );
  NOR2X1 U4172 ( .A(n4677), .B(n4473), .Y(n4675) );
  MXI2X1 U4173 ( .A(n4678), .B(n4679), .S0(randd[25]), .Y(n4673) );
  OAI21X1 U4174 ( .A0(IDtReg[25]), .A1(n4478), .B0(n4479), .Y(n4679) );
  NOR2X1 U4175 ( .A(n4680), .B(n4478), .Y(n4678) );
  MXI2X1 U4176 ( .A(n4681), .B(n4682), .S0(rand_in[25]), .Y(n4672) );
  OAI22X1 U4177 ( .A0(IDtReg[25]), .A1(n4487), .B0(IDstReg[25]), .B1(n4488), 
        .Y(n4682) );
  OAI2B2X1 U4178 ( .A1N(IDstReg[25]), .A0(n4488), .B0(n4680), .B1(n4487), .Y(
        n4681) );
  CLKINVX1 U4179 ( .A(IDtReg[25]), .Y(n4680) );
  MXI2X1 U4180 ( .A(n4683), .B(n4684), .S0(rand_in[57]), .Y(n4671) );
  OAI22X1 U4181 ( .A0(IDtReg[57]), .A1(n4483), .B0(IDstReg[57]), .B1(n4484), 
        .Y(n4684) );
  OAI2B2X1 U4182 ( .A1N(IDstReg[57]), .A0(n4484), .B0(n4677), .B1(n4483), .Y(
        n4683) );
  CLKINVX1 U4183 ( .A(IDtReg[57]), .Y(n4677) );
  NAND4X1 U4184 ( .A(n4685), .B(n4686), .C(n4687), .D(n4688), .Y(
        Inst_AEAD_key[24]) );
  MXI2X1 U4185 ( .A(n4689), .B(n4690), .S0(randd[56]), .Y(n4688) );
  OAI21X1 U4186 ( .A0(IDtReg[56]), .A1(n4473), .B0(n4474), .Y(n4690) );
  NOR2X1 U4187 ( .A(n4691), .B(n4473), .Y(n4689) );
  MXI2X1 U4188 ( .A(n4692), .B(n4693), .S0(randd[24]), .Y(n4687) );
  OAI21X1 U4189 ( .A0(IDtReg[24]), .A1(n4478), .B0(n4479), .Y(n4693) );
  NOR2X1 U4190 ( .A(n4694), .B(n4478), .Y(n4692) );
  MXI2X1 U4191 ( .A(n4695), .B(n4696), .S0(rand_in[24]), .Y(n4686) );
  OAI22X1 U4192 ( .A0(IDtReg[24]), .A1(n4487), .B0(IDstReg[24]), .B1(n4488), 
        .Y(n4696) );
  OAI2B2X1 U4193 ( .A1N(IDstReg[24]), .A0(n4488), .B0(n4694), .B1(n4487), .Y(
        n4695) );
  CLKINVX1 U4194 ( .A(IDtReg[24]), .Y(n4694) );
  MXI2X1 U4195 ( .A(n4697), .B(n4698), .S0(rand_in[56]), .Y(n4685) );
  OAI22X1 U4196 ( .A0(IDtReg[56]), .A1(n4483), .B0(IDstReg[56]), .B1(n4484), 
        .Y(n4698) );
  OAI2B2X1 U4197 ( .A1N(IDstReg[56]), .A0(n4484), .B0(n4691), .B1(n4483), .Y(
        n4697) );
  CLKINVX1 U4198 ( .A(IDtReg[56]), .Y(n4691) );
  NAND4X1 U4199 ( .A(n4699), .B(n4700), .C(n4701), .D(n4702), .Y(
        Inst_AEAD_key[23]) );
  MXI2X1 U4200 ( .A(n4703), .B(n4704), .S0(randd[55]), .Y(n4702) );
  OAI21X1 U4201 ( .A0(IDtReg[55]), .A1(n4473), .B0(n4474), .Y(n4704) );
  NOR2X1 U4202 ( .A(n4705), .B(n4473), .Y(n4703) );
  MXI2X1 U4203 ( .A(n4706), .B(n4707), .S0(randd[23]), .Y(n4701) );
  OAI21X1 U4204 ( .A0(IDtReg[23]), .A1(n4478), .B0(n4479), .Y(n4707) );
  NOR2X1 U4205 ( .A(n4708), .B(n4478), .Y(n4706) );
  MXI2X1 U4206 ( .A(n4709), .B(n4710), .S0(rand_in[23]), .Y(n4700) );
  OAI22X1 U4207 ( .A0(IDtReg[23]), .A1(n4487), .B0(IDstReg[23]), .B1(n4488), 
        .Y(n4710) );
  OAI2B2X1 U4208 ( .A1N(IDstReg[23]), .A0(n4488), .B0(n4708), .B1(n4487), .Y(
        n4709) );
  CLKINVX1 U4209 ( .A(IDtReg[23]), .Y(n4708) );
  MXI2X1 U4210 ( .A(n4711), .B(n4712), .S0(rand_in[55]), .Y(n4699) );
  OAI22X1 U4211 ( .A0(IDtReg[55]), .A1(n4483), .B0(IDstReg[55]), .B1(n4484), 
        .Y(n4712) );
  OAI2B2X1 U4212 ( .A1N(IDstReg[55]), .A0(n4484), .B0(n4705), .B1(n4483), .Y(
        n4711) );
  CLKINVX1 U4213 ( .A(IDtReg[55]), .Y(n4705) );
  NAND4X1 U4214 ( .A(n4713), .B(n4714), .C(n4715), .D(n4716), .Y(
        Inst_AEAD_key[22]) );
  MXI2X1 U4215 ( .A(n4717), .B(n4718), .S0(randd[54]), .Y(n4716) );
  OAI21X1 U4216 ( .A0(IDtReg[54]), .A1(n4473), .B0(n4474), .Y(n4718) );
  NOR2X1 U4217 ( .A(n4719), .B(n4473), .Y(n4717) );
  MXI2X1 U4218 ( .A(n4720), .B(n4721), .S0(randd[22]), .Y(n4715) );
  OAI21X1 U4219 ( .A0(IDtReg[22]), .A1(n4478), .B0(n4479), .Y(n4721) );
  NOR2X1 U4220 ( .A(n4722), .B(n4478), .Y(n4720) );
  MXI2X1 U4221 ( .A(n4723), .B(n4724), .S0(rand_in[22]), .Y(n4714) );
  OAI22X1 U4222 ( .A0(IDtReg[22]), .A1(n4487), .B0(IDstReg[22]), .B1(n4488), 
        .Y(n4724) );
  OAI2B2X1 U4223 ( .A1N(IDstReg[22]), .A0(n4488), .B0(n4722), .B1(n4487), .Y(
        n4723) );
  CLKINVX1 U4224 ( .A(IDtReg[22]), .Y(n4722) );
  MXI2X1 U4225 ( .A(n4725), .B(n4726), .S0(rand_in[54]), .Y(n4713) );
  OAI22X1 U4226 ( .A0(IDtReg[54]), .A1(n4483), .B0(IDstReg[54]), .B1(n4484), 
        .Y(n4726) );
  OAI2B2X1 U4227 ( .A1N(IDstReg[54]), .A0(n4484), .B0(n4719), .B1(n4483), .Y(
        n4725) );
  CLKINVX1 U4228 ( .A(IDtReg[54]), .Y(n4719) );
  NAND4X1 U4229 ( .A(n4727), .B(n4728), .C(n4729), .D(n4730), .Y(
        Inst_AEAD_key[21]) );
  MXI2X1 U4230 ( .A(n4731), .B(n4732), .S0(randd[53]), .Y(n4730) );
  OAI21X1 U4231 ( .A0(IDtReg[53]), .A1(n4473), .B0(n4474), .Y(n4732) );
  NOR2X1 U4232 ( .A(n4733), .B(n4473), .Y(n4731) );
  MXI2X1 U4233 ( .A(n4734), .B(n4735), .S0(randd[21]), .Y(n4729) );
  OAI21X1 U4234 ( .A0(IDtReg[21]), .A1(n4478), .B0(n4479), .Y(n4735) );
  NOR2X1 U4235 ( .A(n4736), .B(n4478), .Y(n4734) );
  MXI2X1 U4236 ( .A(n4737), .B(n4738), .S0(rand_in[21]), .Y(n4728) );
  OAI22X1 U4237 ( .A0(IDtReg[21]), .A1(n4487), .B0(IDstReg[21]), .B1(n4488), 
        .Y(n4738) );
  OAI2B2X1 U4238 ( .A1N(IDstReg[21]), .A0(n4488), .B0(n4736), .B1(n4487), .Y(
        n4737) );
  CLKINVX1 U4239 ( .A(IDtReg[21]), .Y(n4736) );
  MXI2X1 U4240 ( .A(n4739), .B(n4740), .S0(rand_in[53]), .Y(n4727) );
  OAI22X1 U4241 ( .A0(IDtReg[53]), .A1(n4483), .B0(IDstReg[53]), .B1(n4484), 
        .Y(n4740) );
  OAI2B2X1 U4242 ( .A1N(IDstReg[53]), .A0(n4484), .B0(n4733), .B1(n4483), .Y(
        n4739) );
  CLKINVX1 U4243 ( .A(IDtReg[53]), .Y(n4733) );
  NAND4X1 U4244 ( .A(n4741), .B(n4742), .C(n4743), .D(n4744), .Y(
        Inst_AEAD_key[20]) );
  MXI2X1 U4245 ( .A(n4745), .B(n4746), .S0(randd[52]), .Y(n4744) );
  OAI21X1 U4246 ( .A0(IDtReg[52]), .A1(n4473), .B0(n4474), .Y(n4746) );
  NOR2X1 U4247 ( .A(n4747), .B(n4473), .Y(n4745) );
  MXI2X1 U4248 ( .A(n4748), .B(n4749), .S0(randd[20]), .Y(n4743) );
  OAI21X1 U4249 ( .A0(IDtReg[20]), .A1(n4478), .B0(n4479), .Y(n4749) );
  NOR2X1 U4250 ( .A(n4750), .B(n4478), .Y(n4748) );
  MXI2X1 U4251 ( .A(n4751), .B(n4752), .S0(rand_in[20]), .Y(n4742) );
  OAI22X1 U4252 ( .A0(IDtReg[20]), .A1(n4487), .B0(IDstReg[20]), .B1(n4488), 
        .Y(n4752) );
  OAI2B2X1 U4253 ( .A1N(IDstReg[20]), .A0(n4488), .B0(n4750), .B1(n4487), .Y(
        n4751) );
  CLKINVX1 U4254 ( .A(IDtReg[20]), .Y(n4750) );
  MXI2X1 U4255 ( .A(n4753), .B(n4754), .S0(rand_in[52]), .Y(n4741) );
  OAI22X1 U4256 ( .A0(IDtReg[52]), .A1(n4483), .B0(IDstReg[52]), .B1(n4484), 
        .Y(n4754) );
  OAI2B2X1 U4257 ( .A1N(IDstReg[52]), .A0(n4484), .B0(n4747), .B1(n4483), .Y(
        n4753) );
  CLKINVX1 U4258 ( .A(IDtReg[52]), .Y(n4747) );
  NAND4X1 U4259 ( .A(n4755), .B(n4756), .C(n4757), .D(n4758), .Y(
        Inst_AEAD_key[1]) );
  MXI2X1 U4260 ( .A(n4759), .B(n4760), .S0(randd[33]), .Y(n4758) );
  OAI21X1 U4261 ( .A0(IDtReg[33]), .A1(n4473), .B0(n4474), .Y(n4760) );
  NOR2X1 U4262 ( .A(n4761), .B(n4473), .Y(n4759) );
  MXI2X1 U4263 ( .A(n4762), .B(n4763), .S0(randd[1]), .Y(n4757) );
  OAI21X1 U4264 ( .A0(IDtReg[1]), .A1(n4478), .B0(n4479), .Y(n4763) );
  NOR2X1 U4265 ( .A(n4764), .B(n4478), .Y(n4762) );
  MXI2X1 U4266 ( .A(n4765), .B(n4766), .S0(rand_in[1]), .Y(n4756) );
  OAI22X1 U4267 ( .A0(IDtReg[1]), .A1(n4487), .B0(IDstReg[1]), .B1(n4488), .Y(
        n4766) );
  OAI2B2X1 U4268 ( .A1N(IDstReg[1]), .A0(n4488), .B0(n4764), .B1(n4487), .Y(
        n4765) );
  CLKINVX1 U4269 ( .A(IDtReg[1]), .Y(n4764) );
  MXI2X1 U4270 ( .A(n4767), .B(n4768), .S0(rand_in[33]), .Y(n4755) );
  OAI22X1 U4271 ( .A0(IDtReg[33]), .A1(n4483), .B0(IDstReg[33]), .B1(n4484), 
        .Y(n4768) );
  OAI2B2X1 U4272 ( .A1N(IDstReg[33]), .A0(n4484), .B0(n4761), .B1(n4483), .Y(
        n4767) );
  CLKINVX1 U4273 ( .A(IDtReg[33]), .Y(n4761) );
  NAND4X1 U4274 ( .A(n4769), .B(n4770), .C(n4771), .D(n4772), .Y(
        Inst_AEAD_key[19]) );
  MXI2X1 U4275 ( .A(n4773), .B(n4774), .S0(randd[51]), .Y(n4772) );
  OAI21X1 U4276 ( .A0(IDtReg[51]), .A1(n4473), .B0(n4474), .Y(n4774) );
  NOR2X1 U4277 ( .A(n4775), .B(n4473), .Y(n4773) );
  MXI2X1 U4278 ( .A(n4776), .B(n4777), .S0(randd[19]), .Y(n4771) );
  OAI21X1 U4279 ( .A0(IDtReg[19]), .A1(n4478), .B0(n4479), .Y(n4777) );
  NOR2X1 U4280 ( .A(n4778), .B(n4478), .Y(n4776) );
  MXI2X1 U4281 ( .A(n4779), .B(n4780), .S0(rand_in[19]), .Y(n4770) );
  OAI22X1 U4282 ( .A0(IDtReg[19]), .A1(n4487), .B0(IDstReg[19]), .B1(n4488), 
        .Y(n4780) );
  OAI2B2X1 U4283 ( .A1N(IDstReg[19]), .A0(n4488), .B0(n4778), .B1(n4487), .Y(
        n4779) );
  CLKINVX1 U4284 ( .A(IDtReg[19]), .Y(n4778) );
  MXI2X1 U4285 ( .A(n4781), .B(n4782), .S0(rand_in[51]), .Y(n4769) );
  OAI22X1 U4286 ( .A0(IDtReg[51]), .A1(n4483), .B0(IDstReg[51]), .B1(n4484), 
        .Y(n4782) );
  OAI2B2X1 U4287 ( .A1N(IDstReg[51]), .A0(n4484), .B0(n4775), .B1(n4483), .Y(
        n4781) );
  CLKINVX1 U4288 ( .A(IDtReg[51]), .Y(n4775) );
  NAND4X1 U4289 ( .A(n4783), .B(n4784), .C(n4785), .D(n4786), .Y(
        Inst_AEAD_key[18]) );
  MXI2X1 U4290 ( .A(n4787), .B(n4788), .S0(randd[50]), .Y(n4786) );
  OAI21X1 U4291 ( .A0(IDtReg[50]), .A1(n4473), .B0(n4474), .Y(n4788) );
  NOR2X1 U4292 ( .A(n4789), .B(n4473), .Y(n4787) );
  MXI2X1 U4293 ( .A(n4790), .B(n4791), .S0(randd[18]), .Y(n4785) );
  OAI21X1 U4294 ( .A0(IDtReg[18]), .A1(n4478), .B0(n4479), .Y(n4791) );
  NOR2X1 U4295 ( .A(n4792), .B(n4478), .Y(n4790) );
  MXI2X1 U4296 ( .A(n4793), .B(n4794), .S0(rand_in[18]), .Y(n4784) );
  OAI22X1 U4297 ( .A0(IDtReg[18]), .A1(n4487), .B0(IDstReg[18]), .B1(n4488), 
        .Y(n4794) );
  OAI2B2X1 U4298 ( .A1N(IDstReg[18]), .A0(n4488), .B0(n4792), .B1(n4487), .Y(
        n4793) );
  CLKINVX1 U4299 ( .A(IDtReg[18]), .Y(n4792) );
  MXI2X1 U4300 ( .A(n4795), .B(n4796), .S0(rand_in[50]), .Y(n4783) );
  OAI22X1 U4301 ( .A0(IDtReg[50]), .A1(n4483), .B0(IDstReg[50]), .B1(n4484), 
        .Y(n4796) );
  OAI2B2X1 U4302 ( .A1N(IDstReg[50]), .A0(n4484), .B0(n4789), .B1(n4483), .Y(
        n4795) );
  CLKINVX1 U4303 ( .A(IDtReg[50]), .Y(n4789) );
  NAND4X1 U4304 ( .A(n4797), .B(n4798), .C(n4799), .D(n4800), .Y(
        Inst_AEAD_key[17]) );
  MXI2X1 U4305 ( .A(n4801), .B(n4802), .S0(randd[49]), .Y(n4800) );
  OAI21X1 U4306 ( .A0(IDtReg[49]), .A1(n4473), .B0(n4474), .Y(n4802) );
  NOR2X1 U4307 ( .A(n4803), .B(n4473), .Y(n4801) );
  MXI2X1 U4308 ( .A(n4804), .B(n4805), .S0(randd[17]), .Y(n4799) );
  OAI21X1 U4309 ( .A0(IDtReg[17]), .A1(n4478), .B0(n4479), .Y(n4805) );
  NOR2X1 U4310 ( .A(n4806), .B(n4478), .Y(n4804) );
  MXI2X1 U4311 ( .A(n4807), .B(n4808), .S0(rand_in[17]), .Y(n4798) );
  OAI22X1 U4312 ( .A0(IDtReg[17]), .A1(n4487), .B0(IDstReg[17]), .B1(n4488), 
        .Y(n4808) );
  OAI2B2X1 U4313 ( .A1N(IDstReg[17]), .A0(n4488), .B0(n4806), .B1(n4487), .Y(
        n4807) );
  CLKINVX1 U4314 ( .A(IDtReg[17]), .Y(n4806) );
  MXI2X1 U4315 ( .A(n4809), .B(n4810), .S0(rand_in[49]), .Y(n4797) );
  OAI22X1 U4316 ( .A0(IDtReg[49]), .A1(n4483), .B0(IDstReg[49]), .B1(n4484), 
        .Y(n4810) );
  OAI2B2X1 U4317 ( .A1N(IDstReg[49]), .A0(n4484), .B0(n4803), .B1(n4483), .Y(
        n4809) );
  CLKINVX1 U4318 ( .A(IDtReg[49]), .Y(n4803) );
  NAND4X1 U4319 ( .A(n4811), .B(n4812), .C(n4813), .D(n4814), .Y(
        Inst_AEAD_key[16]) );
  MXI2X1 U4320 ( .A(n4815), .B(n4816), .S0(randd[48]), .Y(n4814) );
  OAI21X1 U4321 ( .A0(IDtReg[48]), .A1(n4473), .B0(n4474), .Y(n4816) );
  NOR2X1 U4322 ( .A(n4817), .B(n4473), .Y(n4815) );
  MXI2X1 U4323 ( .A(n4818), .B(n4819), .S0(randd[16]), .Y(n4813) );
  OAI21X1 U4324 ( .A0(IDtReg[16]), .A1(n4478), .B0(n4479), .Y(n4819) );
  NOR2X1 U4325 ( .A(n4820), .B(n4478), .Y(n4818) );
  MXI2X1 U4326 ( .A(n4821), .B(n4822), .S0(rand_in[16]), .Y(n4812) );
  OAI22X1 U4327 ( .A0(IDtReg[16]), .A1(n4487), .B0(IDstReg[16]), .B1(n4488), 
        .Y(n4822) );
  OAI2B2X1 U4328 ( .A1N(IDstReg[16]), .A0(n4488), .B0(n4820), .B1(n4487), .Y(
        n4821) );
  CLKINVX1 U4329 ( .A(IDtReg[16]), .Y(n4820) );
  MXI2X1 U4330 ( .A(n4823), .B(n4824), .S0(rand_in[48]), .Y(n4811) );
  OAI22X1 U4331 ( .A0(IDtReg[48]), .A1(n4483), .B0(IDstReg[48]), .B1(n4484), 
        .Y(n4824) );
  OAI2B2X1 U4332 ( .A1N(IDstReg[48]), .A0(n4484), .B0(n4817), .B1(n4483), .Y(
        n4823) );
  CLKINVX1 U4333 ( .A(IDtReg[48]), .Y(n4817) );
  NAND4X1 U4334 ( .A(n4825), .B(n4826), .C(n4827), .D(n4828), .Y(
        Inst_AEAD_key[15]) );
  MXI2X1 U4335 ( .A(n4829), .B(n4830), .S0(randd[47]), .Y(n4828) );
  OAI21X1 U4336 ( .A0(IDtReg[47]), .A1(n4473), .B0(n4474), .Y(n4830) );
  NOR2X1 U4337 ( .A(n4831), .B(n4473), .Y(n4829) );
  MXI2X1 U4338 ( .A(n4832), .B(n4833), .S0(randd[15]), .Y(n4827) );
  OAI21X1 U4339 ( .A0(IDtReg[15]), .A1(n4478), .B0(n4479), .Y(n4833) );
  NOR2X1 U4340 ( .A(n4834), .B(n4478), .Y(n4832) );
  MXI2X1 U4341 ( .A(n4835), .B(n4836), .S0(rand_in[15]), .Y(n4826) );
  OAI22X1 U4342 ( .A0(IDtReg[15]), .A1(n4487), .B0(IDstReg[15]), .B1(n4488), 
        .Y(n4836) );
  OAI2B2X1 U4343 ( .A1N(IDstReg[15]), .A0(n4488), .B0(n4834), .B1(n4487), .Y(
        n4835) );
  CLKINVX1 U4344 ( .A(IDtReg[15]), .Y(n4834) );
  MXI2X1 U4345 ( .A(n4837), .B(n4838), .S0(rand_in[47]), .Y(n4825) );
  OAI22X1 U4346 ( .A0(IDtReg[47]), .A1(n4483), .B0(IDstReg[47]), .B1(n4484), 
        .Y(n4838) );
  OAI2B2X1 U4347 ( .A1N(IDstReg[47]), .A0(n4484), .B0(n4831), .B1(n4483), .Y(
        n4837) );
  CLKINVX1 U4348 ( .A(IDtReg[47]), .Y(n4831) );
  NAND4X1 U4349 ( .A(n4839), .B(n4840), .C(n4841), .D(n4842), .Y(
        Inst_AEAD_key[14]) );
  MXI2X1 U4350 ( .A(n4843), .B(n4844), .S0(randd[46]), .Y(n4842) );
  OAI21X1 U4351 ( .A0(IDtReg[46]), .A1(n4473), .B0(n4474), .Y(n4844) );
  NOR2X1 U4352 ( .A(n4845), .B(n4473), .Y(n4843) );
  MXI2X1 U4353 ( .A(n4846), .B(n4847), .S0(randd[14]), .Y(n4841) );
  OAI21X1 U4354 ( .A0(IDtReg[14]), .A1(n4478), .B0(n4479), .Y(n4847) );
  NOR2X1 U4355 ( .A(n4848), .B(n4478), .Y(n4846) );
  MXI2X1 U4356 ( .A(n4849), .B(n4850), .S0(rand_in[14]), .Y(n4840) );
  OAI22X1 U4357 ( .A0(IDtReg[14]), .A1(n4487), .B0(IDstReg[14]), .B1(n4488), 
        .Y(n4850) );
  OAI2B2X1 U4358 ( .A1N(IDstReg[14]), .A0(n4488), .B0(n4848), .B1(n4487), .Y(
        n4849) );
  CLKINVX1 U4359 ( .A(IDtReg[14]), .Y(n4848) );
  MXI2X1 U4360 ( .A(n4851), .B(n4852), .S0(rand_in[46]), .Y(n4839) );
  OAI22X1 U4361 ( .A0(IDtReg[46]), .A1(n4483), .B0(IDstReg[46]), .B1(n4484), 
        .Y(n4852) );
  OAI2B2X1 U4362 ( .A1N(IDstReg[46]), .A0(n4484), .B0(n4845), .B1(n4483), .Y(
        n4851) );
  CLKINVX1 U4363 ( .A(IDtReg[46]), .Y(n4845) );
  NAND4X1 U4364 ( .A(n4853), .B(n4854), .C(n4855), .D(n4856), .Y(
        Inst_AEAD_key[13]) );
  MXI2X1 U4365 ( .A(n4857), .B(n4858), .S0(randd[45]), .Y(n4856) );
  OAI21X1 U4366 ( .A0(IDtReg[45]), .A1(n4473), .B0(n4474), .Y(n4858) );
  NOR2X1 U4367 ( .A(n4859), .B(n4473), .Y(n4857) );
  MXI2X1 U4368 ( .A(n4860), .B(n4861), .S0(randd[13]), .Y(n4855) );
  OAI21X1 U4369 ( .A0(IDtReg[13]), .A1(n4478), .B0(n4479), .Y(n4861) );
  NOR2X1 U4370 ( .A(n4862), .B(n4478), .Y(n4860) );
  MXI2X1 U4371 ( .A(n4863), .B(n4864), .S0(rand_in[13]), .Y(n4854) );
  OAI22X1 U4372 ( .A0(IDtReg[13]), .A1(n4487), .B0(IDstReg[13]), .B1(n4488), 
        .Y(n4864) );
  OAI2B2X1 U4373 ( .A1N(IDstReg[13]), .A0(n4488), .B0(n4862), .B1(n4487), .Y(
        n4863) );
  CLKINVX1 U4374 ( .A(IDtReg[13]), .Y(n4862) );
  MXI2X1 U4375 ( .A(n4865), .B(n4866), .S0(rand_in[45]), .Y(n4853) );
  OAI22X1 U4376 ( .A0(IDtReg[45]), .A1(n4483), .B0(IDstReg[45]), .B1(n4484), 
        .Y(n4866) );
  OAI2B2X1 U4377 ( .A1N(IDstReg[45]), .A0(n4484), .B0(n4859), .B1(n4483), .Y(
        n4865) );
  CLKINVX1 U4378 ( .A(IDtReg[45]), .Y(n4859) );
  NAND4X1 U4379 ( .A(n4867), .B(n4868), .C(n4869), .D(n4870), .Y(
        Inst_AEAD_key[12]) );
  MXI2X1 U4380 ( .A(n4871), .B(n4872), .S0(randd[44]), .Y(n4870) );
  OAI21X1 U4381 ( .A0(IDtReg[44]), .A1(n4473), .B0(n4474), .Y(n4872) );
  NOR2X1 U4382 ( .A(n4873), .B(n4473), .Y(n4871) );
  MXI2X1 U4383 ( .A(n4874), .B(n4875), .S0(randd[12]), .Y(n4869) );
  OAI21X1 U4384 ( .A0(IDtReg[12]), .A1(n4478), .B0(n4479), .Y(n4875) );
  NOR2X1 U4385 ( .A(n4876), .B(n4478), .Y(n4874) );
  MXI2X1 U4386 ( .A(n4877), .B(n4878), .S0(rand_in[12]), .Y(n4868) );
  OAI22X1 U4387 ( .A0(IDtReg[12]), .A1(n4487), .B0(IDstReg[12]), .B1(n4488), 
        .Y(n4878) );
  OAI2B2X1 U4388 ( .A1N(IDstReg[12]), .A0(n4488), .B0(n4876), .B1(n4487), .Y(
        n4877) );
  CLKINVX1 U4389 ( .A(IDtReg[12]), .Y(n4876) );
  MXI2X1 U4390 ( .A(n4879), .B(n4880), .S0(rand_in[44]), .Y(n4867) );
  OAI22X1 U4391 ( .A0(IDtReg[44]), .A1(n4483), .B0(IDstReg[44]), .B1(n4484), 
        .Y(n4880) );
  OAI2B2X1 U4392 ( .A1N(IDstReg[44]), .A0(n4484), .B0(n4873), .B1(n4483), .Y(
        n4879) );
  CLKINVX1 U4393 ( .A(IDtReg[44]), .Y(n4873) );
  NAND4X1 U4394 ( .A(n4881), .B(n4882), .C(n4883), .D(n4884), .Y(
        Inst_AEAD_key[11]) );
  MXI2X1 U4395 ( .A(n4885), .B(n4886), .S0(randd[43]), .Y(n4884) );
  OAI21X1 U4396 ( .A0(IDtReg[43]), .A1(n4473), .B0(n4474), .Y(n4886) );
  NOR2X1 U4397 ( .A(n4887), .B(n4473), .Y(n4885) );
  MXI2X1 U4398 ( .A(n4888), .B(n4889), .S0(randd[11]), .Y(n4883) );
  OAI21X1 U4399 ( .A0(IDtReg[11]), .A1(n4478), .B0(n4479), .Y(n4889) );
  NOR2X1 U4400 ( .A(n4890), .B(n4478), .Y(n4888) );
  MXI2X1 U4401 ( .A(n4891), .B(n4892), .S0(rand_in[11]), .Y(n4882) );
  OAI22X1 U4402 ( .A0(IDtReg[11]), .A1(n4487), .B0(IDstReg[11]), .B1(n4488), 
        .Y(n4892) );
  OAI2B2X1 U4403 ( .A1N(IDstReg[11]), .A0(n4488), .B0(n4890), .B1(n4487), .Y(
        n4891) );
  CLKINVX1 U4404 ( .A(IDtReg[11]), .Y(n4890) );
  MXI2X1 U4405 ( .A(n4893), .B(n4894), .S0(rand_in[43]), .Y(n4881) );
  OAI22X1 U4406 ( .A0(IDtReg[43]), .A1(n4483), .B0(IDstReg[43]), .B1(n4484), 
        .Y(n4894) );
  OAI2B2X1 U4407 ( .A1N(IDstReg[43]), .A0(n4484), .B0(n4887), .B1(n4483), .Y(
        n4893) );
  CLKINVX1 U4408 ( .A(IDtReg[43]), .Y(n4887) );
  NAND4X1 U4409 ( .A(n4895), .B(n4896), .C(n4897), .D(n4898), .Y(
        Inst_AEAD_key[10]) );
  MXI2X1 U4410 ( .A(n4899), .B(n4900), .S0(randd[42]), .Y(n4898) );
  OAI21X1 U4411 ( .A0(IDtReg[42]), .A1(n4473), .B0(n4474), .Y(n4900) );
  NOR2X1 U4412 ( .A(n4901), .B(n4473), .Y(n4899) );
  MXI2X1 U4413 ( .A(n4902), .B(n4903), .S0(randd[10]), .Y(n4897) );
  OAI21X1 U4414 ( .A0(IDtReg[10]), .A1(n4478), .B0(n4479), .Y(n4903) );
  NOR2X1 U4415 ( .A(n4904), .B(n4478), .Y(n4902) );
  MXI2X1 U4416 ( .A(n4905), .B(n4906), .S0(rand_in[10]), .Y(n4896) );
  OAI22X1 U4417 ( .A0(IDtReg[10]), .A1(n4487), .B0(IDstReg[10]), .B1(n4488), 
        .Y(n4906) );
  OAI2B2X1 U4418 ( .A1N(IDstReg[10]), .A0(n4488), .B0(n4904), .B1(n4487), .Y(
        n4905) );
  CLKINVX1 U4419 ( .A(IDtReg[10]), .Y(n4904) );
  MXI2X1 U4420 ( .A(n4907), .B(n4908), .S0(rand_in[42]), .Y(n4895) );
  OAI22X1 U4421 ( .A0(IDtReg[42]), .A1(n4483), .B0(IDstReg[42]), .B1(n4484), 
        .Y(n4908) );
  OAI2B2X1 U4422 ( .A1N(IDstReg[42]), .A0(n4484), .B0(n4901), .B1(n4483), .Y(
        n4907) );
  CLKINVX1 U4423 ( .A(IDtReg[42]), .Y(n4901) );
  NAND4X1 U4424 ( .A(n4909), .B(n4910), .C(n4911), .D(n4912), .Y(
        Inst_AEAD_key[0]) );
  MXI2X1 U4425 ( .A(n4913), .B(n4914), .S0(randd[32]), .Y(n4912) );
  OAI21X1 U4426 ( .A0(IDtReg[32]), .A1(n4473), .B0(n4474), .Y(n4914) );
  NOR2X1 U4427 ( .A(n4916), .B(n4473), .Y(n4913) );
  MXI2X1 U4428 ( .A(n4918), .B(n4919), .S0(randd[0]), .Y(n4911) );
  OAI21X1 U4429 ( .A0(IDtReg[0]), .A1(n4478), .B0(n4479), .Y(n4919) );
  NOR2X1 U4430 ( .A(n4921), .B(n4478), .Y(n4918) );
  CLKINVX1 U4431 ( .A(MuxSel2), .Y(n4917) );
  MXI2X1 U4432 ( .A(n4922), .B(n4923), .S0(rand_in[0]), .Y(n4910) );
  OAI22X1 U4433 ( .A0(IDtReg[0]), .A1(n4487), .B0(IDstReg[0]), .B1(n4488), .Y(
        n4923) );
  OAI2B2X1 U4434 ( .A1N(IDstReg[0]), .A0(n4488), .B0(n4921), .B1(n4487), .Y(
        n4922) );
  CLKNAND2X2 U4435 ( .A(DtSel), .B(n4924), .Y(n4487) );
  CLKINVX1 U4436 ( .A(IDtReg[0]), .Y(n4921) );
  CLKNAND2X2 U4437 ( .A(n4924), .B(n4925), .Y(n4488) );
  NOR2X1 U4438 ( .A(n4915), .B(MuxSel1[0]), .Y(n4924) );
  MXI2X1 U4439 ( .A(n4926), .B(n4927), .S0(rand_in[32]), .Y(n4909) );
  OAI22X1 U4440 ( .A0(IDtReg[32]), .A1(n4483), .B0(IDstReg[32]), .B1(n4484), 
        .Y(n4927) );
  OAI2B2X1 U4441 ( .A1N(IDstReg[32]), .A0(n4484), .B0(n4916), .B1(n4483), .Y(
        n4926) );
  CLKNAND2X2 U4442 ( .A(n4928), .B(DtSel), .Y(n4483) );
  CLKINVX1 U4443 ( .A(IDtReg[32]), .Y(n4916) );
  CLKNAND2X2 U4444 ( .A(n4928), .B(n4925), .Y(n4484) );
  CLKINVX1 U4445 ( .A(DtSel), .Y(n4925) );
  NOR2X1 U4446 ( .A(n4915), .B(n4920), .Y(n4928) );
  CLKINVX1 U4447 ( .A(MuxSel1[0]), .Y(n4920) );
  CLKINVX1 U4448 ( .A(MuxSel1[1]), .Y(n4915) );
  OAI221X1 U4449 ( .A0(n1773), .A1(n442), .B0(n2899), .B1(n2900), .C0(n4344), 
        .Y(Inst_AEAD_bdo_valid) );
  NAND3XL U4450 ( .A(Inst_AEAD_bdo_ready), .B(n4370), .C(
        Inst_AEAD_u_cc_u_cc_ctrl_n52), .Y(n4344) );
  NOR2X1 U4451 ( .A(n1608), .B(n879), .Y(n4370) );
  CLKINVX1 U4452 ( .A(Inst_AEAD_u_cc_sel_tag[1]), .Y(n1608) );
  CLKNAND2X2 U4453 ( .A(n1776), .B(n4380), .Y(n2900) );
  CLKINVX1 U4454 ( .A(n4381), .Y(n1776) );
  CLKNAND2X2 U4455 ( .A(n4347), .B(n4364), .Y(n4381) );
  AOI2BB1X1 U4456 ( .A0N(n4929), .A1N(n4930), .B0(n4371), .Y(n4364) );
  CLKINVX1 U4457 ( .A(Inst_AEAD_bdi_valid), .Y(n4371) );
  NAND3XL U4458 ( .A(Inst_AEAD_bdi_size[2]), .B(Inst_AEAD_bdi_size[1]), .C(
        Inst_AEAD_bdi_size[3]), .Y(n4930) );
  NAND3BX1 U4459 ( .AN(Inst_AEAD_bdo_ready), .B(n4380), .C(
        Inst_AEAD_bdi_size[0]), .Y(n4929) );
  CLKNAND2X2 U4460 ( .A(n1564), .B(Inst_AEAD_u_input_n358), .Y(n4380) );
  NOR2X1 U4461 ( .A(n879), .B(Inst_AEAD_u_cc_sel_tag[1]), .Y(n4347) );
  NOR4X1 U4462 ( .A(Inst_AEAD_bdi_size[0]), .B(Inst_AEAD_bdi_size[1]), .C(
        Inst_AEAD_bdi_size[2]), .D(Inst_AEAD_bdi_size[3]), .Y(n2899) );
  NAND3XL U4463 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .B(n4355), .C(
        Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .Y(n1773) );
  OAI222X1 U4464 ( .A0(n2023), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2749), .C0(n1855), .C1(n4932), .Y(Inst_AEAD_bdo[9]) );
  XNOR2X1 U4465 ( .A(n4933), .B(n1251), .Y(n1855) );
  NAND2BX1 U4466 ( .AN(n1137), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4933) );
  XNOR2X1 U4467 ( .A(Inst_AEAD_u_input_n313), .B(n1506), .Y(n2749) );
  XNOR2X1 U4468 ( .A(n4934), .B(n1314), .Y(n2023) );
  NAND2BX1 U4469 ( .AN(n1139), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4934) );
  OAI222X1 U4470 ( .A0(n2030), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2759), .C0(n1919), .C1(n4932), .Y(Inst_AEAD_bdo[8]) );
  XNOR2X1 U4471 ( .A(n4935), .B(n1250), .Y(n1919) );
  NAND2BX1 U4472 ( .AN(n1141), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4935) );
  XNOR2X1 U4473 ( .A(Inst_AEAD_u_input_n314), .B(n1505), .Y(n2759) );
  XNOR2X1 U4474 ( .A(n4936), .B(n1313), .Y(n2030) );
  NAND2BX1 U4475 ( .AN(n1143), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4936) );
  OAI222X1 U4476 ( .A0(n2037), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2776), .C0(n1974), .C1(n4932), .Y(Inst_AEAD_bdo[7]) );
  XNOR2X1 U4477 ( .A(n4937), .B(n1249), .Y(n1974) );
  NAND2BX1 U4478 ( .AN(n1145), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4937) );
  XNOR2X1 U4479 ( .A(n1976), .B(n1504), .Y(n2776) );
  CLKINVX1 U4480 ( .A(Inst_AEAD_bdi[7]), .Y(n1976) );
  XNOR2X1 U4481 ( .A(n4938), .B(n1312), .Y(n2037) );
  NAND2BX1 U4482 ( .AN(n1147), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4938) );
  OAI222X1 U4483 ( .A0(n2045), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2796), .C0(n2053), .C1(n4932), .Y(Inst_AEAD_bdo[6]) );
  XNOR2X1 U4484 ( .A(n4939), .B(n1248), .Y(n2053) );
  NAND2BX1 U4485 ( .AN(n1149), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4939) );
  XNOR2X1 U4486 ( .A(Inst_AEAD_u_input_n315), .B(n1503), .Y(n2796) );
  XNOR2X1 U4487 ( .A(n4940), .B(n1311), .Y(n2045) );
  NAND2BX1 U4488 ( .AN(n1151), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4940) );
  OAI222X1 U4489 ( .A0(n4176), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n4941), .C0(n2106), .C1(n4932), .Y(Inst_AEAD_bdo[63]) );
  XNOR2X1 U4490 ( .A(n4942), .B(n1305), .Y(n2106) );
  NAND2BX1 U4491 ( .AN(n1050), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4942) );
  XNOR2X1 U4492 ( .A(n1560), .B(n1600), .Y(n4941) );
  XNOR2X1 U4493 ( .A(n4943), .B(n1368), .Y(n4176) );
  NAND2BX1 U4494 ( .AN(n1052), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4943) );
  OAI222X1 U4495 ( .A0(n4181), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2296), .C0(n2111), .C1(n4932), .Y(Inst_AEAD_bdo[62]) );
  XNOR2X1 U4496 ( .A(n4944), .B(n1304), .Y(n2111) );
  NAND2BX1 U4497 ( .AN(n1054), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4944) );
  XNOR2X1 U4498 ( .A(n1559), .B(n1568), .Y(n2296) );
  XNOR2X1 U4499 ( .A(n4945), .B(n1367), .Y(n4181) );
  NAND2BX1 U4500 ( .AN(n1056), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4945) );
  OAI222X1 U4501 ( .A0(n4186), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2303), .C0(n2117), .C1(n4932), .Y(Inst_AEAD_bdo[61]) );
  XNOR2X1 U4502 ( .A(n4946), .B(n1303), .Y(n2117) );
  NAND2BX1 U4503 ( .AN(n1058), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4946) );
  XNOR2X1 U4504 ( .A(n1558), .B(n1569), .Y(n2303) );
  XNOR2X1 U4505 ( .A(n4947), .B(n1366), .Y(n4186) );
  NAND2BX1 U4506 ( .AN(n1060), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4947) );
  OAI222X1 U4507 ( .A0(n4191), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2309), .C0(n2123), .C1(n4932), .Y(Inst_AEAD_bdo[60]) );
  XNOR2X1 U4508 ( .A(n4948), .B(n1302), .Y(n2123) );
  NAND2BX1 U4509 ( .AN(n1062), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4948) );
  XNOR2X1 U4510 ( .A(n1557), .B(n1570), .Y(n2309) );
  XNOR2X1 U4511 ( .A(n4949), .B(n1365), .Y(n4191) );
  NAND2BX1 U4512 ( .AN(n1064), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4949) );
  OAI222X1 U4513 ( .A0(n2059), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2812), .C0(n2129), .C1(n4932), .Y(Inst_AEAD_bdo[5]) );
  XNOR2X1 U4514 ( .A(n4950), .B(n1247), .Y(n2129) );
  NAND2BX1 U4515 ( .AN(n1153), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4950) );
  XNOR2X1 U4516 ( .A(Inst_AEAD_u_input_n316), .B(n1502), .Y(n2812) );
  XNOR2X1 U4517 ( .A(n4951), .B(n1310), .Y(n2059) );
  NAND2BX1 U4518 ( .AN(n1155), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4951) );
  OAI222X1 U4519 ( .A0(n4196), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2315), .C0(n2134), .C1(n4932), .Y(Inst_AEAD_bdo[59]) );
  XNOR2X1 U4520 ( .A(n4952), .B(n1301), .Y(n2134) );
  NAND2BX1 U4521 ( .AN(n1066), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4952) );
  XNOR2X1 U4522 ( .A(n1556), .B(n1571), .Y(n2315) );
  XNOR2X1 U4523 ( .A(n4953), .B(n1364), .Y(n4196) );
  NAND2BX1 U4524 ( .AN(n1068), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4953) );
  OAI222X1 U4525 ( .A0(n4201), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2321), .C0(n2140), .C1(n4932), .Y(Inst_AEAD_bdo[58]) );
  XNOR2X1 U4526 ( .A(n4954), .B(n1300), .Y(n2140) );
  NAND2BX1 U4527 ( .AN(n1070), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4954) );
  XNOR2X1 U4528 ( .A(n1555), .B(n1572), .Y(n2321) );
  XNOR2X1 U4529 ( .A(n4955), .B(n1363), .Y(n4201) );
  NAND2BX1 U4530 ( .AN(n1072), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4955) );
  OAI222X1 U4531 ( .A0(n4207), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2327), .C0(n2146), .C1(n4932), .Y(Inst_AEAD_bdo[57]) );
  XNOR2X1 U4532 ( .A(n4956), .B(n1299), .Y(n2146) );
  NAND2BX1 U4533 ( .AN(n1074), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4956) );
  XNOR2X1 U4534 ( .A(n1554), .B(n1573), .Y(n2327) );
  XNOR2X1 U4535 ( .A(n4957), .B(n1362), .Y(n4207) );
  NAND2BX1 U4536 ( .AN(n1076), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4957) );
  OAI222X1 U4537 ( .A0(n4213), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2333), .C0(n2152), .C1(n4932), .Y(Inst_AEAD_bdo[56]) );
  XNOR2X1 U4538 ( .A(n4958), .B(n1298), .Y(n2152) );
  NAND2BX1 U4539 ( .AN(n1078), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4958) );
  XNOR2X1 U4540 ( .A(n1553), .B(n1574), .Y(n2333) );
  XNOR2X1 U4541 ( .A(n4959), .B(n1361), .Y(n4213) );
  NAND2BX1 U4542 ( .AN(n1080), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4959) );
  OAI222X1 U4543 ( .A0(n4221), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2341), .C0(n2157), .C1(n4932), .Y(Inst_AEAD_bdo[55]) );
  XNOR2X1 U4544 ( .A(n4960), .B(n1297), .Y(n2157) );
  NAND2BX1 U4545 ( .AN(n1082), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4960) );
  XNOR2X1 U4546 ( .A(n1552), .B(n1601), .Y(n2341) );
  XNOR2X1 U4547 ( .A(n4961), .B(n1360), .Y(n4221) );
  NAND2BX1 U4548 ( .AN(n1084), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4961) );
  OAI222X1 U4549 ( .A0(n4226), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n4962), .C0(n2162), .C1(n4932), .Y(Inst_AEAD_bdo[54]) );
  XNOR2X1 U4550 ( .A(n4963), .B(n1296), .Y(n2162) );
  NAND2BX1 U4551 ( .AN(n1086), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4963) );
  XNOR2X1 U4552 ( .A(n1551), .B(n1575), .Y(n4962) );
  XNOR2X1 U4553 ( .A(n4964), .B(n1359), .Y(n4226) );
  NAND2BX1 U4554 ( .AN(n1088), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4964) );
  OAI222X1 U4555 ( .A0(n4233), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2361), .C0(n2167), .C1(n4932), .Y(Inst_AEAD_bdo[53]) );
  XNOR2X1 U4556 ( .A(n4965), .B(n1295), .Y(n2167) );
  NAND2BX1 U4557 ( .AN(n1090), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4965) );
  XNOR2X1 U4558 ( .A(n1550), .B(n1576), .Y(n2361) );
  XNOR2X1 U4559 ( .A(n4966), .B(n1358), .Y(n4233) );
  NAND2BX1 U4560 ( .AN(n1092), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4966) );
  OAI222X1 U4561 ( .A0(n4238), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2366), .C0(n2172), .C1(n4932), .Y(Inst_AEAD_bdo[52]) );
  XNOR2X1 U4562 ( .A(n4967), .B(n1294), .Y(n2172) );
  NAND2BX1 U4563 ( .AN(n1094), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4967) );
  XNOR2X1 U4564 ( .A(n1549), .B(n1577), .Y(n2366) );
  XNOR2X1 U4565 ( .A(n4968), .B(n1357), .Y(n4238) );
  NAND2BX1 U4566 ( .AN(n1096), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4968) );
  OAI222X1 U4567 ( .A0(n4243), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2371), .C0(n2177), .C1(n4932), .Y(Inst_AEAD_bdo[51]) );
  XNOR2X1 U4568 ( .A(n4969), .B(n1293), .Y(n2177) );
  NAND2BX1 U4569 ( .AN(n1098), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4969) );
  XNOR2X1 U4570 ( .A(n1548), .B(n1578), .Y(n2371) );
  XNOR2X1 U4571 ( .A(n4970), .B(n1356), .Y(n4243) );
  NAND2BX1 U4572 ( .AN(n1100), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4970) );
  OAI222X1 U4573 ( .A0(n4247), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2376), .C0(n2182), .C1(n4932), .Y(Inst_AEAD_bdo[50]) );
  XNOR2X1 U4574 ( .A(n4971), .B(n1292), .Y(n2182) );
  NAND2BX1 U4575 ( .AN(n1102), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4971) );
  XNOR2X1 U4576 ( .A(n1547), .B(n1579), .Y(n2376) );
  XNOR2X1 U4577 ( .A(n4972), .B(n1355), .Y(n4247) );
  NAND2BX1 U4578 ( .AN(n1104), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4972) );
  OAI222X1 U4579 ( .A0(n2067), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2828), .C0(n2186), .C1(n4932), .Y(Inst_AEAD_bdo[4]) );
  XNOR2X1 U4580 ( .A(n4973), .B(n1246), .Y(n2186) );
  NAND2BX1 U4581 ( .AN(n1157), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4973) );
  XNOR2X1 U4582 ( .A(Inst_AEAD_u_input_n317), .B(n1501), .Y(n2828) );
  XNOR2X1 U4583 ( .A(n4974), .B(n1309), .Y(n2067) );
  NAND2BX1 U4584 ( .AN(n1159), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4974) );
  OAI222X1 U4585 ( .A0(n4251), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2381), .C0(n2191), .C1(n4932), .Y(Inst_AEAD_bdo[49]) );
  XNOR2X1 U4586 ( .A(n4975), .B(n1291), .Y(n2191) );
  NAND2BX1 U4587 ( .AN(n1106), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4975) );
  XNOR2X1 U4588 ( .A(n1546), .B(n1580), .Y(n2381) );
  XNOR2X1 U4589 ( .A(n4976), .B(n1354), .Y(n4251) );
  NAND2BX1 U4590 ( .AN(n1108), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4976) );
  OAI222X1 U4591 ( .A0(n4255), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2386), .C0(n2195), .C1(n4932), .Y(Inst_AEAD_bdo[48]) );
  XNOR2X1 U4592 ( .A(n4977), .B(n1290), .Y(n2195) );
  NAND2BX1 U4593 ( .AN(n1110), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4977) );
  XNOR2X1 U4594 ( .A(n1545), .B(n1581), .Y(n2386) );
  XNOR2X1 U4595 ( .A(n4978), .B(n1353), .Y(n4255) );
  NAND2BX1 U4596 ( .AN(n1112), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4978) );
  OAI222X1 U4597 ( .A0(n4259), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2391), .C0(n2199), .C1(n4932), .Y(Inst_AEAD_bdo[47]) );
  XNOR2X1 U4598 ( .A(n4979), .B(n1289), .Y(n2199) );
  NAND2BX1 U4599 ( .AN(n1114), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4979) );
  XNOR2X1 U4600 ( .A(n1544), .B(n1602), .Y(n2391) );
  XNOR2X1 U4601 ( .A(n4980), .B(n1352), .Y(n4259) );
  NAND2BX1 U4602 ( .AN(n1116), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4980) );
  OAI222X1 U4603 ( .A0(n4263), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2398), .C0(n2203), .C1(n4932), .Y(Inst_AEAD_bdo[46]) );
  XNOR2X1 U4604 ( .A(n4981), .B(n1288), .Y(n2203) );
  NAND2BX1 U4605 ( .AN(n1118), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4981) );
  XNOR2X1 U4606 ( .A(n1543), .B(n1582), .Y(n2398) );
  XNOR2X1 U4607 ( .A(n4982), .B(n1351), .Y(n4263) );
  NAND2BX1 U4608 ( .AN(n1120), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4982) );
  OAI222X1 U4609 ( .A0(n4270), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2403), .C0(n2207), .C1(n4932), .Y(Inst_AEAD_bdo[45]) );
  XNOR2X1 U4610 ( .A(n4983), .B(n1287), .Y(n2207) );
  NAND2BX1 U4611 ( .AN(n1122), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4983) );
  XNOR2X1 U4612 ( .A(n1542), .B(n1583), .Y(n2403) );
  XNOR2X1 U4613 ( .A(n4984), .B(n1350), .Y(n4270) );
  NAND2BX1 U4614 ( .AN(n1124), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4984) );
  OAI222X1 U4615 ( .A0(n4275), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2408), .C0(n2211), .C1(n4932), .Y(Inst_AEAD_bdo[44]) );
  XNOR2X1 U4616 ( .A(n4985), .B(n1286), .Y(n2211) );
  NAND2BX1 U4617 ( .AN(n1126), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4985) );
  XNOR2X1 U4618 ( .A(n1541), .B(n1584), .Y(n2408) );
  XNOR2X1 U4619 ( .A(n4986), .B(n1349), .Y(n4275) );
  NAND2BX1 U4620 ( .AN(n1128), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4986) );
  OAI222X1 U4621 ( .A0(n4280), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n4987), .C0(n2216), .C1(n4932), .Y(Inst_AEAD_bdo[43]) );
  XNOR2X1 U4622 ( .A(n4988), .B(n1285), .Y(n2216) );
  NAND2BX1 U4623 ( .AN(n1130), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4988) );
  XNOR2X1 U4624 ( .A(n1540), .B(n1585), .Y(n4987) );
  XNOR2X1 U4625 ( .A(n4989), .B(n1348), .Y(n4280) );
  NAND2BX1 U4626 ( .AN(n1132), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4989) );
  OAI222X1 U4627 ( .A0(n4285), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n4990), .C0(n2223), .C1(n4932), .Y(Inst_AEAD_bdo[42]) );
  XNOR2X1 U4628 ( .A(n4991), .B(n1284), .Y(n2223) );
  NAND2BX1 U4629 ( .AN(n1134), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4991) );
  XNOR2X1 U4630 ( .A(n1539), .B(n1586), .Y(n4990) );
  XNOR2X1 U4631 ( .A(n4992), .B(n1347), .Y(n4285) );
  NAND2BX1 U4632 ( .AN(n1136), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4992) );
  OAI222X1 U4633 ( .A0(n4291), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2440), .C0(n2230), .C1(n4932), .Y(Inst_AEAD_bdo[41]) );
  XNOR2X1 U4634 ( .A(n4993), .B(n1283), .Y(n2230) );
  NAND2BX1 U4635 ( .AN(n1138), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4993) );
  XNOR2X1 U4636 ( .A(n1538), .B(n1587), .Y(n2440) );
  XNOR2X1 U4637 ( .A(n4994), .B(n1346), .Y(n4291) );
  NAND2BX1 U4638 ( .AN(n1140), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4994) );
  OAI222X1 U4639 ( .A0(n4297), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2444), .C0(n2237), .C1(n4932), .Y(Inst_AEAD_bdo[40]) );
  XNOR2X1 U4640 ( .A(n4995), .B(n1282), .Y(n2237) );
  NAND2BX1 U4641 ( .AN(n1142), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4995) );
  XNOR2X1 U4642 ( .A(n1537), .B(n1588), .Y(n2444) );
  XNOR2X1 U4643 ( .A(n4996), .B(n1345), .Y(n4297) );
  NAND2BX1 U4644 ( .AN(n1144), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4996) );
  OAI222X1 U4645 ( .A0(n2075), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2851), .C0(n2243), .C1(n4932), .Y(Inst_AEAD_bdo[3]) );
  XNOR2X1 U4646 ( .A(n4997), .B(n1245), .Y(n2243) );
  NAND2BX1 U4647 ( .AN(n1161), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4997) );
  XNOR2X1 U4648 ( .A(Inst_AEAD_u_input_n318), .B(n1500), .Y(n2851) );
  XNOR2X1 U4649 ( .A(n4998), .B(n1308), .Y(n2075) );
  NAND2BX1 U4650 ( .AN(n1163), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4998) );
  OAI222X1 U4651 ( .A0(n4303), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2448), .C0(n2247), .C1(n4932), .Y(Inst_AEAD_bdo[39]) );
  XNOR2X1 U4652 ( .A(n4999), .B(n1281), .Y(n2247) );
  NAND2BX1 U4653 ( .AN(n1146), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n4999) );
  XNOR2X1 U4654 ( .A(n1536), .B(n1603), .Y(n2448) );
  XNOR2X1 U4655 ( .A(n5000), .B(n1344), .Y(n4303) );
  NAND2BX1 U4656 ( .AN(n1148), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5000) );
  OAI222X1 U4657 ( .A0(n4309), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2454), .C0(n2252), .C1(n4932), .Y(Inst_AEAD_bdo[38]) );
  XNOR2X1 U4658 ( .A(n5001), .B(n1280), .Y(n2252) );
  NAND2BX1 U4659 ( .AN(n1150), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5001) );
  XNOR2X1 U4660 ( .A(n1535), .B(n1589), .Y(n2454) );
  XNOR2X1 U4661 ( .A(n5002), .B(n1343), .Y(n4309) );
  NAND2BX1 U4662 ( .AN(n1152), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5002) );
  OAI222X1 U4663 ( .A0(n4315), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2458), .C0(n2257), .C1(n4932), .Y(Inst_AEAD_bdo[37]) );
  XNOR2X1 U4664 ( .A(n5003), .B(n1279), .Y(n2257) );
  NAND2BX1 U4665 ( .AN(n1154), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5003) );
  XNOR2X1 U4666 ( .A(n1534), .B(n1590), .Y(n2458) );
  XNOR2X1 U4667 ( .A(n5004), .B(n1342), .Y(n4315) );
  NAND2BX1 U4668 ( .AN(n1156), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5004) );
  OAI222X1 U4669 ( .A0(n4321), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2462), .C0(n2262), .C1(n4932), .Y(Inst_AEAD_bdo[36]) );
  XNOR2X1 U4670 ( .A(n5005), .B(n1278), .Y(n2262) );
  NAND2BX1 U4671 ( .AN(n1158), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5005) );
  XNOR2X1 U4672 ( .A(n1533), .B(n1591), .Y(n2462) );
  XNOR2X1 U4673 ( .A(n5006), .B(n1341), .Y(n4321) );
  NAND2BX1 U4674 ( .AN(n1160), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5006) );
  OAI222X1 U4675 ( .A0(n1862), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2466), .C0(n2265), .C1(n4932), .Y(Inst_AEAD_bdo[35]) );
  XNOR2X1 U4676 ( .A(n5007), .B(n1277), .Y(n2265) );
  NAND2BX1 U4677 ( .AN(n1162), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5007) );
  XNOR2X1 U4678 ( .A(n1532), .B(n1592), .Y(n2466) );
  XNOR2X1 U4679 ( .A(n5008), .B(n1340), .Y(n1862) );
  NAND2BX1 U4680 ( .AN(n1164), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5008) );
  OAI222X1 U4681 ( .A0(n1868), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n5009), .C0(n2268), .C1(n4932), .Y(Inst_AEAD_bdo[34]) );
  XNOR2X1 U4682 ( .A(n5010), .B(n1276), .Y(n2268) );
  NAND2BX1 U4683 ( .AN(n1166), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5010) );
  XNOR2X1 U4684 ( .A(n1531), .B(n1593), .Y(n5009) );
  XNOR2X1 U4685 ( .A(n5011), .B(n1339), .Y(n1868) );
  NAND2BX1 U4686 ( .AN(n1168), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5011) );
  OAI222X1 U4687 ( .A0(n1874), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n5012), .C0(n2271), .C1(n4932), .Y(Inst_AEAD_bdo[33]) );
  XNOR2X1 U4688 ( .A(n5013), .B(n1275), .Y(n2271) );
  NAND2BX1 U4689 ( .AN(n1170), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5013) );
  XNOR2X1 U4690 ( .A(n1530), .B(n1594), .Y(n5012) );
  XNOR2X1 U4691 ( .A(n5014), .B(n1338), .Y(n1874) );
  NAND2BX1 U4692 ( .AN(n1172), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5014) );
  OAI222X1 U4693 ( .A0(n1880), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2505), .C0(n2276), .C1(n4932), .Y(Inst_AEAD_bdo[32]) );
  XNOR2X1 U4694 ( .A(n5015), .B(n1274), .Y(n2276) );
  NAND2BX1 U4695 ( .AN(n1174), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5015) );
  XNOR2X1 U4696 ( .A(n1529), .B(n1595), .Y(n2505) );
  XNOR2X1 U4697 ( .A(n5016), .B(n1337), .Y(n1880) );
  NAND2BX1 U4698 ( .AN(n1176), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5016) );
  OAI222X1 U4699 ( .A0(n1886), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2515), .C0(n2281), .C1(n4932), .Y(Inst_AEAD_bdo[31]) );
  XNOR2X1 U4700 ( .A(n5017), .B(n1273), .Y(n2281) );
  NAND2BX1 U4701 ( .AN(n1049), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5017) );
  XNOR2X1 U4702 ( .A(Inst_AEAD_u_input_n303), .B(n1528), .Y(n2515) );
  XNOR2X1 U4703 ( .A(n5018), .B(n1336), .Y(n1886) );
  NAND2BX1 U4704 ( .AN(n1051), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5018) );
  OAI222X1 U4705 ( .A0(n1892), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2525), .C0(n2355), .C1(n4932), .Y(Inst_AEAD_bdo[30]) );
  XNOR2X1 U4706 ( .A(n5019), .B(n1272), .Y(n2355) );
  NAND2BX1 U4707 ( .AN(n1053), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5019) );
  XNOR2X1 U4708 ( .A(Inst_AEAD_u_input_n304), .B(n1527), .Y(n2525) );
  XNOR2X1 U4709 ( .A(n5020), .B(n1335), .Y(n1892) );
  NAND2BX1 U4710 ( .AN(n1055), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5020) );
  OAI222X1 U4711 ( .A0(n2083), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2866), .C0(n2411), .C1(n4932), .Y(Inst_AEAD_bdo[2]) );
  XNOR2X1 U4712 ( .A(n5021), .B(n1244), .Y(n2411) );
  NAND2BX1 U4713 ( .AN(n1165), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5021) );
  XNOR2X1 U4714 ( .A(Inst_AEAD_u_input_n319), .B(n1499), .Y(n2866) );
  XNOR2X1 U4715 ( .A(n5022), .B(n1307), .Y(n2083) );
  NAND2BX1 U4716 ( .AN(n1167), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5022) );
  OAI222X1 U4717 ( .A0(n1898), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2534), .C0(n2418), .C1(n4932), .Y(Inst_AEAD_bdo[29]) );
  XNOR2X1 U4718 ( .A(n5023), .B(n1271), .Y(n2418) );
  NAND2BX1 U4719 ( .AN(n1057), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5023) );
  XNOR2X1 U4720 ( .A(Inst_AEAD_u_input_n305), .B(n1526), .Y(n2534) );
  XNOR2X1 U4721 ( .A(n5024), .B(n1334), .Y(n1898) );
  NAND2BX1 U4722 ( .AN(n1059), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5024) );
  OAI222X1 U4723 ( .A0(n1904), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2543), .C0(n2486), .C1(n4932), .Y(Inst_AEAD_bdo[28]) );
  XNOR2X1 U4724 ( .A(n5025), .B(n1270), .Y(n2486) );
  NAND2BX1 U4725 ( .AN(n1061), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5025) );
  XNOR2X1 U4726 ( .A(Inst_AEAD_u_input_n306), .B(n1525), .Y(n2543) );
  XNOR2X1 U4727 ( .A(n5026), .B(n1333), .Y(n1904) );
  NAND2BX1 U4728 ( .AN(n1063), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5026) );
  OAI222X1 U4729 ( .A0(n1909), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2552), .C0(n2585), .C1(n4932), .Y(Inst_AEAD_bdo[27]) );
  XNOR2X1 U4730 ( .A(n5027), .B(n1269), .Y(n2585) );
  NAND2BX1 U4731 ( .AN(n1065), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5027) );
  XNOR2X1 U4732 ( .A(n1726), .B(n1524), .Y(n2552) );
  CLKINVX1 U4733 ( .A(Inst_AEAD_bdi[27]), .Y(n1726) );
  XNOR2X1 U4734 ( .A(n5028), .B(n1332), .Y(n1909) );
  NAND2BX1 U4735 ( .AN(n1067), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5028) );
  OAI222X1 U4736 ( .A0(n1914), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2560), .C0(n2694), .C1(n4932), .Y(Inst_AEAD_bdo[26]) );
  XNOR2X1 U4737 ( .A(n5029), .B(n1268), .Y(n2694) );
  NAND2BX1 U4738 ( .AN(n1069), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5029) );
  XNOR2X1 U4739 ( .A(n1725), .B(n1523), .Y(n2560) );
  CLKINVX1 U4740 ( .A(Inst_AEAD_bdi[26]), .Y(n1725) );
  XNOR2X1 U4741 ( .A(n5030), .B(n1331), .Y(n1914) );
  NAND2BX1 U4742 ( .AN(n1071), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5030) );
  OAI222X1 U4743 ( .A0(n1925), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2568), .C0(n2844), .C1(n4932), .Y(Inst_AEAD_bdo[25]) );
  XNOR2X1 U4744 ( .A(n5031), .B(n1267), .Y(n2844) );
  NAND2BX1 U4745 ( .AN(n1073), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5031) );
  XNOR2X1 U4746 ( .A(Inst_AEAD_u_input_n307), .B(n1522), .Y(n2568) );
  XNOR2X1 U4747 ( .A(n5032), .B(n1330), .Y(n1925) );
  NAND2BX1 U4748 ( .AN(n1075), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5032) );
  OAI222X1 U4749 ( .A0(n1929), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2576), .C0(n2956), .C1(n4932), .Y(Inst_AEAD_bdo[24]) );
  XNOR2X1 U4750 ( .A(n5033), .B(n1266), .Y(n2956) );
  NAND2BX1 U4751 ( .AN(n1077), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5033) );
  XNOR2X1 U4752 ( .A(n1722), .B(n1521), .Y(n2576) );
  CLKINVX1 U4753 ( .A(Inst_AEAD_bdi[24]), .Y(n1722) );
  XNOR2X1 U4754 ( .A(n5034), .B(n1329), .Y(n1929) );
  NAND2BX1 U4755 ( .AN(n1079), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5034) );
  OAI222X1 U4756 ( .A0(n1933), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2594), .C0(n3020), .C1(n4932), .Y(Inst_AEAD_bdo[23]) );
  XNOR2X1 U4757 ( .A(n5035), .B(n1265), .Y(n3020) );
  NAND2BX1 U4758 ( .AN(n1081), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5035) );
  XNOR2X1 U4759 ( .A(n2595), .B(n1520), .Y(n2594) );
  CLKINVX1 U4760 ( .A(Inst_AEAD_bdi[23]), .Y(n2595) );
  XNOR2X1 U4761 ( .A(n5036), .B(n1328), .Y(n1933) );
  NAND2BX1 U4762 ( .AN(n1083), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5036) );
  OAI222X1 U4763 ( .A0(n1937), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2605), .C0(n3086), .C1(n4932), .Y(Inst_AEAD_bdo[22]) );
  XNOR2X1 U4764 ( .A(n5037), .B(n1264), .Y(n3086) );
  NAND2BX1 U4765 ( .AN(n1085), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5037) );
  XNOR2X1 U4766 ( .A(n1721), .B(n1519), .Y(n2605) );
  CLKINVX1 U4767 ( .A(Inst_AEAD_bdi[22]), .Y(n1721) );
  XNOR2X1 U4768 ( .A(n5038), .B(n1327), .Y(n1937) );
  NAND2BX1 U4769 ( .AN(n1087), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5038) );
  OAI222X1 U4770 ( .A0(n1941), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2612), .C0(n3211), .C1(n4932), .Y(Inst_AEAD_bdo[21]) );
  XNOR2X1 U4771 ( .A(n5039), .B(n1263), .Y(n3211) );
  NAND2BX1 U4772 ( .AN(n1089), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5039) );
  XNOR2X1 U4773 ( .A(n1720), .B(n1518), .Y(n2612) );
  CLKINVX1 U4774 ( .A(Inst_AEAD_bdi[21]), .Y(n1720) );
  XNOR2X1 U4775 ( .A(n5040), .B(n1326), .Y(n1941) );
  NAND2BX1 U4776 ( .AN(n1091), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5040) );
  OAI222X1 U4777 ( .A0(n1945), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2619), .C0(n3366), .C1(n4932), .Y(Inst_AEAD_bdo[20]) );
  XNOR2X1 U4778 ( .A(n5041), .B(n1262), .Y(n3366) );
  NAND2BX1 U4779 ( .AN(n1093), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5041) );
  XNOR2X1 U4780 ( .A(n1719), .B(n1517), .Y(n2619) );
  CLKINVX1 U4781 ( .A(Inst_AEAD_bdi[20]), .Y(n1719) );
  XNOR2X1 U4782 ( .A(n5042), .B(n1325), .Y(n1945) );
  NAND2BX1 U4783 ( .AN(n1095), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5042) );
  OAI222X1 U4784 ( .A0(n2091), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2881), .C0(n3561), .C1(n4932), .Y(Inst_AEAD_bdo[1]) );
  XNOR2X1 U4785 ( .A(n5043), .B(n1243), .Y(n3561) );
  NAND2BX1 U4786 ( .AN(n1169), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5043) );
  XNOR2X1 U4787 ( .A(Inst_AEAD_u_input_n320), .B(n1498), .Y(n2881) );
  XNOR2X1 U4788 ( .A(n5044), .B(n1306), .Y(n2091) );
  NAND2BX1 U4789 ( .AN(n1171), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5044) );
  OAI222X1 U4790 ( .A0(n1949), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2626), .C0(n3566), .C1(n4932), .Y(Inst_AEAD_bdo[19]) );
  XNOR2X1 U4791 ( .A(n5045), .B(n1261), .Y(n3566) );
  NAND2BX1 U4792 ( .AN(n1097), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5045) );
  XNOR2X1 U4793 ( .A(n1718), .B(n1516), .Y(n2626) );
  CLKINVX1 U4794 ( .A(Inst_AEAD_bdi[19]), .Y(n1718) );
  XNOR2X1 U4795 ( .A(n5046), .B(n1324), .Y(n1949) );
  NAND2BX1 U4796 ( .AN(n1099), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5046) );
  OAI222X1 U4797 ( .A0(n1953), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2633), .C0(n3752), .C1(n4932), .Y(Inst_AEAD_bdo[18]) );
  XNOR2X1 U4798 ( .A(n5047), .B(n1260), .Y(n3752) );
  NAND2BX1 U4799 ( .AN(n1101), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5047) );
  XNOR2X1 U4800 ( .A(n1717), .B(n1515), .Y(n2633) );
  CLKINVX1 U4801 ( .A(Inst_AEAD_bdi[18]), .Y(n1717) );
  XNOR2X1 U4802 ( .A(n5048), .B(n1323), .Y(n1953) );
  NAND2BX1 U4803 ( .AN(n1103), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5048) );
  OAI222X1 U4804 ( .A0(n1960), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2644), .C0(n3818), .C1(n4932), .Y(Inst_AEAD_bdo[17]) );
  XNOR2X1 U4805 ( .A(n5049), .B(n1259), .Y(n3818) );
  NAND2BX1 U4806 ( .AN(n1105), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5049) );
  XNOR2X1 U4807 ( .A(n1716), .B(n1514), .Y(n2644) );
  CLKINVX1 U4808 ( .A(Inst_AEAD_bdi[17]), .Y(n1716) );
  XNOR2X1 U4809 ( .A(n5050), .B(n1322), .Y(n1960) );
  NAND2BX1 U4810 ( .AN(n1107), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5050) );
  OAI222X1 U4811 ( .A0(n1967), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2655), .C0(n3886), .C1(n4932), .Y(Inst_AEAD_bdo[16]) );
  XNOR2X1 U4812 ( .A(n5051), .B(n1258), .Y(n3886) );
  NAND2BX1 U4813 ( .AN(n1109), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5051) );
  XNOR2X1 U4814 ( .A(n1715), .B(n1513), .Y(n2655) );
  CLKINVX1 U4815 ( .A(Inst_AEAD_bdi[16]), .Y(n1715) );
  XNOR2X1 U4816 ( .A(n5052), .B(n1321), .Y(n1967) );
  NAND2BX1 U4817 ( .AN(n1111), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5052) );
  OAI222X1 U4818 ( .A0(n1981), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2668), .C0(n3959), .C1(n4932), .Y(Inst_AEAD_bdo[15]) );
  XNOR2X1 U4819 ( .A(n5053), .B(n1257), .Y(n3959) );
  NAND2BX1 U4820 ( .AN(n1113), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5053) );
  XNOR2X1 U4821 ( .A(n2669), .B(n1512), .Y(n2668) );
  CLKINVX1 U4822 ( .A(Inst_AEAD_bdi[15]), .Y(n2669) );
  XNOR2X1 U4823 ( .A(n5054), .B(n1320), .Y(n1981) );
  NAND2BX1 U4824 ( .AN(n1115), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5054) );
  OAI222X1 U4825 ( .A0(n1988), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2682), .C0(n4024), .C1(n4932), .Y(Inst_AEAD_bdo[14]) );
  XNOR2X1 U4826 ( .A(n5055), .B(n1256), .Y(n4024) );
  NAND2BX1 U4827 ( .AN(n1117), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5055) );
  XNOR2X1 U4828 ( .A(Inst_AEAD_u_input_n308), .B(n1511), .Y(n2682) );
  XNOR2X1 U4829 ( .A(n5056), .B(n1319), .Y(n1988) );
  NAND2BX1 U4830 ( .AN(n1119), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5056) );
  OAI222X1 U4831 ( .A0(n1995), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2702), .C0(n4087), .C1(n4932), .Y(Inst_AEAD_bdo[13]) );
  XNOR2X1 U4832 ( .A(n5057), .B(n1255), .Y(n4087) );
  NAND2BX1 U4833 ( .AN(n1121), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5057) );
  XNOR2X1 U4834 ( .A(Inst_AEAD_u_input_n309), .B(n1510), .Y(n2702) );
  XNOR2X1 U4835 ( .A(n5058), .B(n1318), .Y(n1995) );
  NAND2BX1 U4836 ( .AN(n1123), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5058) );
  OAI222X1 U4837 ( .A0(n2002), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2715), .C0(n4159), .C1(n4932), .Y(Inst_AEAD_bdo[12]) );
  XNOR2X1 U4838 ( .A(n5059), .B(n1254), .Y(n4159) );
  NAND2BX1 U4839 ( .AN(n1125), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5059) );
  XNOR2X1 U4840 ( .A(Inst_AEAD_u_input_n310), .B(n1509), .Y(n2715) );
  XNOR2X1 U4841 ( .A(n5060), .B(n1317), .Y(n2002) );
  NAND2BX1 U4842 ( .AN(n1127), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5060) );
  OAI222X1 U4843 ( .A0(n2009), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2727), .C0(n4218), .C1(n4932), .Y(Inst_AEAD_bdo[11]) );
  XNOR2X1 U4844 ( .A(n5061), .B(n1253), .Y(n4218) );
  NAND2BX1 U4845 ( .AN(n1129), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5061) );
  XNOR2X1 U4846 ( .A(Inst_AEAD_u_input_n311), .B(n1508), .Y(n2727) );
  XNOR2X1 U4847 ( .A(n5062), .B(n1316), .Y(n2009) );
  NAND2BX1 U4848 ( .AN(n1131), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5062) );
  OAI222X1 U4849 ( .A0(n2016), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2738), .C0(n4267), .C1(n4932), .Y(Inst_AEAD_bdo[10]) );
  XNOR2X1 U4850 ( .A(n5063), .B(n1252), .Y(n4267) );
  NAND2BX1 U4851 ( .AN(n1133), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5063) );
  XNOR2X1 U4852 ( .A(Inst_AEAD_u_input_n312), .B(n1507), .Y(n2738) );
  XNOR2X1 U4853 ( .A(n5064), .B(n1315), .Y(n2016) );
  NAND2BX1 U4854 ( .AN(n1135), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5064) );
  OAI222X1 U4855 ( .A0(n2099), .A1(n4931), .B0(Inst_AEAD_u_cc_sel_tag[1]), 
        .B1(n2898), .C0(n4327), .C1(n4932), .Y(Inst_AEAD_bdo[0]) );
  CLKNAND2X2 U4856 ( .A(Inst_AEAD_u_cc_sel_tag[0]), .B(
        Inst_AEAD_u_cc_sel_tag[1]), .Y(n4932) );
  XNOR2X1 U4857 ( .A(n5065), .B(n5066), .Y(n4327) );
  NOR2BX1 U4858 ( .AN(Inst_AEAD_u_cc_sel_key_lo), .B(n1173), .Y(n5066) );
  XNOR2X1 U4859 ( .A(n1242), .B(n4377), .Y(n5065) );
  NOR4BX1 U4860 ( .AN(Inst_AEAD_u_input_n358), .B(n879), .C(
        Inst_AEAD_u_cc_u_cc_ctrl_is_init_dat), .D(n1564), .Y(n4377) );
  CLKINVX1 U4861 ( .A(n2334), .Y(n1854) );
  NOR3X1 U4862 ( .A(n4355), .B(Inst_AEAD_u_cc_u_cc_ctrl_state_1_), .C(n4352), 
        .Y(n2334) );
  CLKINVX1 U4863 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_2_), .Y(n4352) );
  CLKINVX1 U4864 ( .A(Inst_AEAD_u_cc_u_cc_ctrl_state_0_), .Y(n4355) );
  XNOR2X1 U4865 ( .A(Inst_AEAD_u_input_n321), .B(n1497), .Y(n2898) );
  XNOR2X1 U4866 ( .A(n5067), .B(n1241), .Y(n2099) );
  NAND2BX1 U4867 ( .AN(n1175), .B(Inst_AEAD_u_cc_sel_key_lo), .Y(n5067) );
endmodule


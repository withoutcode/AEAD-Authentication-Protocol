
module Skinny_Imp ( clk, rst, en_c, ld_rec, IDt, IDst, DtSel, rand_in, MuxSel2, 
        a_data, enc, dec, gen_tag, Input1, Input2, N, K1, K2, Block_Size, 
        Output1, Output2, Tag1, Tag2, done );
  input [63:0] IDt;
  input [63:0] IDst;
  input [63:0] rand_in;
  input [127:0] Input1;
  input [127:0] Input2;
  input [95:0] N;
  input [127:0] K1;
  input [127:0] K2;
  input [3:0] Block_Size;
  output [127:0] Output1;
  output [127:0] Output2;
  output [127:0] Tag1;
  output [127:0] Tag2;
  input clk, rst, en_c, ld_rec, DtSel, MuxSel2, a_data, enc, dec, gen_tag;
  output done;
  wire   Inst_forkAE_LFSRInst_n63, Inst_forkAE_LFSRInst_n62,
         Inst_forkAE_LFSRInst_n61, Inst_forkAE_LFSRInst_n52,
         Inst_forkAE_LFSRInst_n51, Inst_forkAE_CipherInst_LAST,
         Inst_forkAE_CipherInst_TK1_DEC_0_, Inst_forkAE_CipherInst_TK1_DEC_1_,
         Inst_forkAE_CipherInst_TK1_DEC_2_, Inst_forkAE_CipherInst_TK1_DEC_3_,
         Inst_forkAE_CipherInst_TK1_DEC_4_, Inst_forkAE_CipherInst_TK1_DEC_5_,
         Inst_forkAE_CipherInst_TK1_DEC_6_, Inst_forkAE_CipherInst_TK1_DEC_7_,
         Inst_forkAE_CipherInst_TK1_DEC_48_,
         Inst_forkAE_CipherInst_TK1_DEC_49_,
         Inst_forkAE_CipherInst_TK1_DEC_51_,
         Inst_forkAE_CipherInst_TK1_DEC_52_,
         Inst_forkAE_CipherInst_TK1_DEC_53_,
         Inst_forkAE_CipherInst_TK1_DEC_54_,
         Inst_forkAE_CipherInst_TK1_DEC_55_,
         Inst_forkAE_CipherInst_TK1_DEC_56_,
         Inst_forkAE_CipherInst_TK1_DEC_57_,
         Inst_forkAE_CipherInst_TK1_DEC_58_,
         Inst_forkAE_CipherInst_TK1_DEC_59_,
         Inst_forkAE_CipherInst_TK1_DEC_60_,
         Inst_forkAE_CipherInst_TK1_DEC_61_,
         Inst_forkAE_CipherInst_TK1_DEC_62_, Inst_forkAE_ControlInst_n33,
         Inst_forkAE_ControlInst_n32, Inst_forkAE_ControlInst_n31,
         Inst_forkAE_ControlInst_encdec_started,
         Inst_forkAE_ControlInst_fsm_state_0_,
         Inst_forkAE_ControlInst_fsm_state_1_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_0_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_1_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_2_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_3_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_4_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_5_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_6_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_7_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_8_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_9_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_10_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_11_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_12_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_13_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_14_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_15_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_16_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_17_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_18_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_19_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_20_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_21_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_22_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_23_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_24_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_25_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_26_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_27_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_28_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_29_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_30_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_31_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_32_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_33_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_34_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_35_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_36_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_37_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_38_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_39_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_40_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_41_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_42_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_43_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_44_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_45_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_46_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_47_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_48_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_49_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_50_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_51_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_52_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_53_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_54_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_55_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_56_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_57_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_58_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_59_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_60_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_61_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_62_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_63_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_64_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_65_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_66_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_67_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_68_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_69_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_70_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_71_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_72_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_73_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_74_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_75_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_76_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_77_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_78_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_79_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_80_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_81_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_82_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_83_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_84_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_85_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_86_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_87_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_88_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_89_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_90_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_91_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_92_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_93_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_94_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_95_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_96_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_97_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_98_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_99_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_100_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_101_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_102_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_103_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_104_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_105_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_106_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_107_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_108_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_109_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_110_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_111_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_112_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_113_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_114_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_115_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_116_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_117_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_118_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_119_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_120_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_121_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_122_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_123_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_124_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_125_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_126_,
         Inst_forkAE_MainPart1_Tag_Reg_Output_127_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_0_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_1_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_2_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_3_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_4_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_5_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_6_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_7_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_8_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_9_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_10_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_11_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_12_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_13_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_14_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_15_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_16_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_17_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_18_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_19_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_20_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_21_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_22_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_23_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_24_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_25_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_26_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_27_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_28_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_29_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_30_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_31_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_32_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_33_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_34_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_35_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_36_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_37_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_38_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_39_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_40_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_41_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_42_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_43_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_44_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_45_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_46_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_47_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_48_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_49_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_50_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_51_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_52_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_53_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_54_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_55_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_56_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_57_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_58_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_59_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_60_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_61_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_62_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_63_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_64_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_65_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_66_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_67_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_68_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_69_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_70_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_71_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_72_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_73_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_74_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_75_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_76_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_77_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_78_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_79_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_80_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_81_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_82_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_83_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_84_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_85_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_86_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_87_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_88_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_89_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_90_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_91_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_92_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_93_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_94_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_95_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_96_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_97_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_98_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_99_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_100_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_101_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_102_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_103_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_104_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_105_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_106_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_107_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_108_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_109_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_110_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_111_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_112_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_113_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_114_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_115_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_116_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_117_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_118_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_119_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_120_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_121_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_122_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_123_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_124_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_125_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_126_,
         Inst_forkAE_MainPart2_Tag_Reg_Output_127_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_0_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_1_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_2_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_3_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_4_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_5_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_6_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_7_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_8_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_9_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_10_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_11_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_12_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_13_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_14_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_15_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_16_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_17_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_18_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_19_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_20_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_21_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_22_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_23_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_24_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_25_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_26_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_27_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_28_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_29_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_30_,
         Inst_forkAE_CipherInst_RF_STATE_EX2_31_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_0_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_1_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_2_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_3_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_4_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_5_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_6_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_7_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_8_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_9_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_10_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_11_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_12_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_13_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_14_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_15_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_16_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_17_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_18_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_19_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_20_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_21_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_22_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_23_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_24_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_25_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_26_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_27_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_28_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_29_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_30_,
         Inst_forkAE_CipherInst_RF_STATE_EX1_31_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_0_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_1_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_2_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_3_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_4_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_5_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_6_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_7_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_8_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_9_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_10_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_11_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_12_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_13_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_14_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_15_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_16_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_17_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_18_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_19_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_20_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_21_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_22_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_23_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_24_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_25_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_26_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_27_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_28_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_29_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_31_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_32_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_33_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_34_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_35_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_36_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_37_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_39_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_40_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_41_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_42_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_43_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_44_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_45_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_47_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_48_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_49_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_50_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_51_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_52_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_53_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_54_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_55_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_56_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_57_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_58_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_59_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_60_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_61_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_62_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_63_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_64_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_65_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_66_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_67_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_68_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_69_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_70_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_71_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_72_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_73_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_74_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_75_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_76_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_77_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_78_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_79_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_80_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_81_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_82_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_83_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_84_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_85_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_86_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_87_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_88_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_89_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_90_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_91_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_92_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_93_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_94_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_95_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_96_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_97_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_98_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_99_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_100_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_101_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_102_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_103_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_104_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_105_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_106_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_107_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_108_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_109_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_110_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_111_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_112_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_113_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_114_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_115_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_116_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_117_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_118_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_119_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_120_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_121_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_122_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_123_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_124_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_125_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_126_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_127_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_0_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_1_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_2_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_3_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_4_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_5_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_6_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_7_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_8_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_9_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_10_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_11_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_12_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_13_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_14_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_15_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_16_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_17_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_18_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_19_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_20_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_21_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_22_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_23_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_24_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_25_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_26_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_27_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_28_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_29_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_30_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_31_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_32_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_33_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_34_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_35_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_36_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_37_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_38_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_39_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_40_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_41_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_42_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_43_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_44_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_45_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_46_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_47_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_48_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_49_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_50_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_51_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_52_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_53_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_54_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_55_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_56_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_57_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_58_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_59_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_60_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_61_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_62_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_63_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_64_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_65_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_66_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_67_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_68_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_69_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_70_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_71_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_72_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_73_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_74_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_75_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_76_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_77_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_78_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_79_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_80_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_81_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_82_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_83_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_84_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_85_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_86_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_87_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_88_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_89_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_90_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_91_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_92_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_93_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_94_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_95_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_96_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_97_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_98_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_99_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_100_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_101_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_102_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_103_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_104_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_105_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_106_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_107_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_108_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_109_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_110_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_111_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_112_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_113_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_114_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_115_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_116_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_117_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_118_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_119_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_120_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_121_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_122_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_123_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_124_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_125_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_126_,
         Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_127_,
         Inst_forkAE_CipherInst_KE_CLK_K, Inst_forkAE_CipherInst_KE_N2,
         Inst_forkAE_CipherInst_CL_n44, Inst_forkAE_CipherInst_CL_n43,
         Inst_forkAE_CipherInst_CL_n34, Inst_forkAE_CipherInst_CL_n27,
         Inst_forkAE_CipherInst_CL_n23, Inst_forkAE_CipherInst_CL_n22,
         Inst_forkAE_CipherInst_CL_STATE_0_, Inst_forkAE_CipherInst_CL_N15,
         Inst_forkAE_CipherInst_CL_N13, Inst_forkAE_CipherInst_CL_COUNTER_0_,
         Inst_forkAE_CipherInst_CL_COUNTER_2_,
         Inst_forkAE_MainPart1_AuthRegInst_n387,
         Inst_forkAE_MainPart1_AuthRegInst_n386,
         Inst_forkAE_MainPart1_AuthRegInst_n385,
         Inst_forkAE_MainPart1_AuthRegInst_n384,
         Inst_forkAE_MainPart1_AuthRegInst_n383,
         Inst_forkAE_MainPart1_AuthRegInst_n382,
         Inst_forkAE_MainPart1_AuthRegInst_n381,
         Inst_forkAE_MainPart1_AuthRegInst_n380,
         Inst_forkAE_MainPart1_AuthRegInst_n379,
         Inst_forkAE_MainPart1_AuthRegInst_n378,
         Inst_forkAE_MainPart1_AuthRegInst_n377,
         Inst_forkAE_MainPart1_AuthRegInst_n376,
         Inst_forkAE_MainPart1_AuthRegInst_n375,
         Inst_forkAE_MainPart1_AuthRegInst_n374,
         Inst_forkAE_MainPart1_AuthRegInst_n373,
         Inst_forkAE_MainPart1_AuthRegInst_n372,
         Inst_forkAE_MainPart1_AuthRegInst_n371,
         Inst_forkAE_MainPart1_AuthRegInst_n370,
         Inst_forkAE_MainPart1_AuthRegInst_n369,
         Inst_forkAE_MainPart1_AuthRegInst_n368,
         Inst_forkAE_MainPart1_AuthRegInst_n367,
         Inst_forkAE_MainPart1_AuthRegInst_n366,
         Inst_forkAE_MainPart1_AuthRegInst_n365,
         Inst_forkAE_MainPart1_AuthRegInst_n364,
         Inst_forkAE_MainPart1_AuthRegInst_n363,
         Inst_forkAE_MainPart1_AuthRegInst_n362,
         Inst_forkAE_MainPart1_AuthRegInst_n361,
         Inst_forkAE_MainPart1_AuthRegInst_n360,
         Inst_forkAE_MainPart1_AuthRegInst_n359,
         Inst_forkAE_MainPart1_AuthRegInst_n358,
         Inst_forkAE_MainPart1_AuthRegInst_n357,
         Inst_forkAE_MainPart1_AuthRegInst_n356,
         Inst_forkAE_MainPart1_AuthRegInst_n355,
         Inst_forkAE_MainPart1_AuthRegInst_n354,
         Inst_forkAE_MainPart1_AuthRegInst_n353,
         Inst_forkAE_MainPart1_AuthRegInst_n352,
         Inst_forkAE_MainPart1_AuthRegInst_n351,
         Inst_forkAE_MainPart1_AuthRegInst_n350,
         Inst_forkAE_MainPart1_AuthRegInst_n349,
         Inst_forkAE_MainPart1_AuthRegInst_n348,
         Inst_forkAE_MainPart1_AuthRegInst_n347,
         Inst_forkAE_MainPart1_AuthRegInst_n346,
         Inst_forkAE_MainPart1_AuthRegInst_n345,
         Inst_forkAE_MainPart1_AuthRegInst_n344,
         Inst_forkAE_MainPart1_AuthRegInst_n343,
         Inst_forkAE_MainPart1_AuthRegInst_n342,
         Inst_forkAE_MainPart1_AuthRegInst_n341,
         Inst_forkAE_MainPart1_AuthRegInst_n340,
         Inst_forkAE_MainPart1_AuthRegInst_n339,
         Inst_forkAE_MainPart1_AuthRegInst_n338,
         Inst_forkAE_MainPart1_AuthRegInst_n337,
         Inst_forkAE_MainPart1_AuthRegInst_n336,
         Inst_forkAE_MainPart1_AuthRegInst_n335,
         Inst_forkAE_MainPart1_AuthRegInst_n334,
         Inst_forkAE_MainPart1_AuthRegInst_n333,
         Inst_forkAE_MainPart1_AuthRegInst_n332,
         Inst_forkAE_MainPart1_AuthRegInst_n331,
         Inst_forkAE_MainPart1_AuthRegInst_n330,
         Inst_forkAE_MainPart1_AuthRegInst_n329,
         Inst_forkAE_MainPart1_AuthRegInst_n328,
         Inst_forkAE_MainPart1_AuthRegInst_n327,
         Inst_forkAE_MainPart1_AuthRegInst_n326,
         Inst_forkAE_MainPart1_AuthRegInst_n325,
         Inst_forkAE_MainPart1_AuthRegInst_n324,
         Inst_forkAE_MainPart1_AuthRegInst_n323,
         Inst_forkAE_MainPart1_AuthRegInst_n322,
         Inst_forkAE_MainPart1_AuthRegInst_n321,
         Inst_forkAE_MainPart1_AuthRegInst_n320,
         Inst_forkAE_MainPart1_AuthRegInst_n319,
         Inst_forkAE_MainPart1_AuthRegInst_n318,
         Inst_forkAE_MainPart1_AuthRegInst_n317,
         Inst_forkAE_MainPart1_AuthRegInst_n316,
         Inst_forkAE_MainPart1_AuthRegInst_n315,
         Inst_forkAE_MainPart1_AuthRegInst_n314,
         Inst_forkAE_MainPart1_AuthRegInst_n313,
         Inst_forkAE_MainPart1_AuthRegInst_n312,
         Inst_forkAE_MainPart1_AuthRegInst_n311,
         Inst_forkAE_MainPart1_AuthRegInst_n310,
         Inst_forkAE_MainPart1_AuthRegInst_n309,
         Inst_forkAE_MainPart1_AuthRegInst_n308,
         Inst_forkAE_MainPart1_AuthRegInst_n307,
         Inst_forkAE_MainPart1_AuthRegInst_n306,
         Inst_forkAE_MainPart1_AuthRegInst_n305,
         Inst_forkAE_MainPart1_AuthRegInst_n304,
         Inst_forkAE_MainPart1_AuthRegInst_n303,
         Inst_forkAE_MainPart1_AuthRegInst_n302,
         Inst_forkAE_MainPart1_AuthRegInst_n301,
         Inst_forkAE_MainPart1_AuthRegInst_n300,
         Inst_forkAE_MainPart1_AuthRegInst_n299,
         Inst_forkAE_MainPart1_AuthRegInst_n298,
         Inst_forkAE_MainPart1_AuthRegInst_n297,
         Inst_forkAE_MainPart1_AuthRegInst_n296,
         Inst_forkAE_MainPart1_AuthRegInst_n295,
         Inst_forkAE_MainPart1_AuthRegInst_n294,
         Inst_forkAE_MainPart1_AuthRegInst_n293,
         Inst_forkAE_MainPart1_AuthRegInst_n292,
         Inst_forkAE_MainPart1_AuthRegInst_n291,
         Inst_forkAE_MainPart1_AuthRegInst_n290,
         Inst_forkAE_MainPart1_AuthRegInst_n289,
         Inst_forkAE_MainPart1_AuthRegInst_n288,
         Inst_forkAE_MainPart1_AuthRegInst_n287,
         Inst_forkAE_MainPart1_AuthRegInst_n286,
         Inst_forkAE_MainPart1_AuthRegInst_n285,
         Inst_forkAE_MainPart1_AuthRegInst_n284,
         Inst_forkAE_MainPart1_AuthRegInst_n283,
         Inst_forkAE_MainPart1_AuthRegInst_n282,
         Inst_forkAE_MainPart1_AuthRegInst_n281,
         Inst_forkAE_MainPart1_AuthRegInst_n280,
         Inst_forkAE_MainPart1_AuthRegInst_n279,
         Inst_forkAE_MainPart1_AuthRegInst_n278,
         Inst_forkAE_MainPart1_AuthRegInst_n277,
         Inst_forkAE_MainPart1_AuthRegInst_n276,
         Inst_forkAE_MainPart1_AuthRegInst_n275,
         Inst_forkAE_MainPart1_AuthRegInst_n274,
         Inst_forkAE_MainPart1_AuthRegInst_n273,
         Inst_forkAE_MainPart1_AuthRegInst_n272,
         Inst_forkAE_MainPart1_AuthRegInst_n271,
         Inst_forkAE_MainPart1_AuthRegInst_n270,
         Inst_forkAE_MainPart1_AuthRegInst_n269,
         Inst_forkAE_MainPart1_AuthRegInst_n268,
         Inst_forkAE_MainPart1_AuthRegInst_n267,
         Inst_forkAE_MainPart1_AuthRegInst_n266,
         Inst_forkAE_MainPart1_AuthRegInst_n265,
         Inst_forkAE_MainPart1_AuthRegInst_n264,
         Inst_forkAE_MainPart1_AuthRegInst_n263,
         Inst_forkAE_MainPart1_AuthRegInst_n262,
         Inst_forkAE_MainPart1_AuthRegInst_n261,
         Inst_forkAE_MainPart1_AuthRegInst_n260,
         Inst_forkAE_CipherInst_RF_RS_EX1_N34,
         Inst_forkAE_CipherInst_RF_RS_EX1_N33,
         Inst_forkAE_CipherInst_RF_RS_EX1_N32,
         Inst_forkAE_CipherInst_RF_RS_EX1_N31,
         Inst_forkAE_CipherInst_RF_RS_EX1_N30,
         Inst_forkAE_CipherInst_RF_RS_EX1_N29,
         Inst_forkAE_CipherInst_RF_RS_EX1_N28,
         Inst_forkAE_CipherInst_RF_RS_EX1_N27,
         Inst_forkAE_CipherInst_RF_RS_EX1_N26,
         Inst_forkAE_CipherInst_RF_RS_EX1_N25,
         Inst_forkAE_CipherInst_RF_RS_EX1_N24,
         Inst_forkAE_CipherInst_RF_RS_EX1_N23,
         Inst_forkAE_CipherInst_RF_RS_EX1_N22,
         Inst_forkAE_CipherInst_RF_RS_EX1_N21,
         Inst_forkAE_CipherInst_RF_RS_EX1_N20,
         Inst_forkAE_CipherInst_RF_RS_EX1_N19,
         Inst_forkAE_CipherInst_RF_RS_EX1_N18,
         Inst_forkAE_CipherInst_RF_RS_EX1_N17,
         Inst_forkAE_CipherInst_RF_RS_EX1_N16,
         Inst_forkAE_CipherInst_RF_RS_EX1_N15,
         Inst_forkAE_CipherInst_RF_RS_EX1_N14,
         Inst_forkAE_CipherInst_RF_RS_EX1_N13,
         Inst_forkAE_CipherInst_RF_RS_EX1_N12,
         Inst_forkAE_CipherInst_RF_RS_EX1_N11,
         Inst_forkAE_CipherInst_RF_RS_EX1_N10,
         Inst_forkAE_CipherInst_RF_RS_EX1_N9,
         Inst_forkAE_CipherInst_RF_RS_EX1_N8,
         Inst_forkAE_CipherInst_RF_RS_EX1_N7,
         Inst_forkAE_CipherInst_RF_RS_EX1_N6,
         Inst_forkAE_CipherInst_RF_RS_EX1_N5,
         Inst_forkAE_CipherInst_RF_RS_EX1_N4,
         Inst_forkAE_CipherInst_RF_RS_EX1_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_0_N3,
         Inst_forkAE_CipherInst_RF_RS_EX2_N34,
         Inst_forkAE_CipherInst_RF_RS_EX2_N33,
         Inst_forkAE_CipherInst_RF_RS_EX2_N32,
         Inst_forkAE_CipherInst_RF_RS_EX2_N31,
         Inst_forkAE_CipherInst_RF_RS_EX2_N30,
         Inst_forkAE_CipherInst_RF_RS_EX2_N29,
         Inst_forkAE_CipherInst_RF_RS_EX2_N28,
         Inst_forkAE_CipherInst_RF_RS_EX2_N27,
         Inst_forkAE_CipherInst_RF_RS_EX2_N26,
         Inst_forkAE_CipherInst_RF_RS_EX2_N25,
         Inst_forkAE_CipherInst_RF_RS_EX2_N24,
         Inst_forkAE_CipherInst_RF_RS_EX2_N23,
         Inst_forkAE_CipherInst_RF_RS_EX2_N22,
         Inst_forkAE_CipherInst_RF_RS_EX2_N21,
         Inst_forkAE_CipherInst_RF_RS_EX2_N20,
         Inst_forkAE_CipherInst_RF_RS_EX2_N19,
         Inst_forkAE_CipherInst_RF_RS_EX2_N18,
         Inst_forkAE_CipherInst_RF_RS_EX2_N17,
         Inst_forkAE_CipherInst_RF_RS_EX2_N16,
         Inst_forkAE_CipherInst_RF_RS_EX2_N15,
         Inst_forkAE_CipherInst_RF_RS_EX2_N14,
         Inst_forkAE_CipherInst_RF_RS_EX2_N13,
         Inst_forkAE_CipherInst_RF_RS_EX2_N12,
         Inst_forkAE_CipherInst_RF_RS_EX2_N11,
         Inst_forkAE_CipherInst_RF_RS_EX2_N10,
         Inst_forkAE_CipherInst_RF_RS_EX2_N9,
         Inst_forkAE_CipherInst_RF_RS_EX2_N8,
         Inst_forkAE_CipherInst_RF_RS_EX2_N7,
         Inst_forkAE_CipherInst_RF_RS_EX2_N6,
         Inst_forkAE_CipherInst_RF_RS_EX2_N5,
         Inst_forkAE_CipherInst_RF_RS_EX2_N4,
         Inst_forkAE_CipherInst_RF_RS_EX2_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_127_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_126_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_125_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_124_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_123_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_122_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_121_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_120_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_119_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_118_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_117_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_116_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_115_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_114_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_113_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_112_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_111_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_110_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_109_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_108_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_107_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_106_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_105_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_104_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_103_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_102_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_101_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_100_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_99_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_98_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_97_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_96_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_95_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_94_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_93_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_92_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_91_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_90_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_89_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_88_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_87_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_86_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_85_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_84_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_83_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_82_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_81_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_80_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_79_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_78_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_77_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_76_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_75_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_74_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_73_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_72_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_71_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_70_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_69_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_68_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_67_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_66_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_65_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_64_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_63_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_62_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_61_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_60_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_59_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_58_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_57_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_56_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_55_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_54_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_53_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_52_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_51_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_50_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_49_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_48_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_47_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_46_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_45_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_44_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_43_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_42_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_41_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_40_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_39_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_38_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_37_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_36_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_35_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_34_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_33_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_32_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_31_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_30_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_29_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_28_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_27_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_26_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_25_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_24_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_23_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_22_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_21_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_20_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_19_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_18_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_17_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_16_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_15_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_14_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_13_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_12_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_11_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_10_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_9_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_8_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_7_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_6_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_5_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_4_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_3_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_2_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_1_N3,
         Inst_forkAE_CipherInst_KE_RS2_2_SFF_0_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_127_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_126_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_125_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_124_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_123_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_122_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_121_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_120_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_119_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_118_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_117_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_116_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_115_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_114_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_113_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_112_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_111_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_110_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_109_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_108_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_107_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_106_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_105_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_104_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_103_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_102_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_101_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_100_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_99_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_98_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_97_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_96_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_95_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_94_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_93_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_92_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_91_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_90_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_89_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_88_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_87_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_86_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_85_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_84_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_83_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_82_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_81_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_80_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_79_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_78_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_77_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_76_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_75_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_74_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_73_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_72_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_71_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_70_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_69_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_68_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_67_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_66_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_65_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_64_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_63_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_62_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_61_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_60_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_59_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_58_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_57_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_56_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_55_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_54_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_53_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_52_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_51_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_50_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_49_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_48_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_47_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_46_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_45_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_44_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_43_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_42_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_41_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_40_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_39_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_38_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_37_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_36_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_35_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_34_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_33_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_32_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_31_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_30_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_29_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_28_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_27_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_26_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_25_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_24_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_23_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_22_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_21_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_20_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_19_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_18_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_17_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_16_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_15_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_14_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_13_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_12_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_11_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_10_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_9_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_8_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_7_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_6_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_5_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_4_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_3_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_2_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_1_N3,
         Inst_forkAE_CipherInst_KE_RS2_1_SFF_0_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_127_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_126_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_125_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_124_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_123_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_122_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_121_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_120_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_119_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_118_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_117_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_116_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_115_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_114_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_113_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_112_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_111_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_110_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_109_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_108_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_107_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_106_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_105_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_104_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_103_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_102_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_101_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_100_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_99_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_98_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_97_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_96_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_95_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_94_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_93_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_92_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_91_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_90_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_89_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_88_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_87_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_86_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_85_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_84_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_83_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_82_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_81_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_80_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_79_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_78_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_77_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_76_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_75_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_74_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_73_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_72_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_71_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_70_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_69_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_68_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_67_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_66_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_65_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_64_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_63_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_62_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_61_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_60_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_59_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_58_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_57_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_56_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_55_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_54_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_53_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_52_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_51_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_50_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_49_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_48_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_47_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_46_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_45_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_44_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_43_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_42_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_41_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_40_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_39_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_38_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_37_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_36_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_35_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_34_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_33_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_32_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_31_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_30_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_29_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_28_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_27_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_26_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_25_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_24_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_23_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_22_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_21_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_20_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_19_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_18_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_17_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_16_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_15_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_14_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_13_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_12_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_11_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_10_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_9_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_8_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_7_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_6_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_5_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_4_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_3_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_2_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_1_N3,
         Inst_forkAE_CipherInst_KE_RS1_SFF_0_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_127_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_126_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_125_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_124_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_123_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_122_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_121_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_120_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_119_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_118_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_117_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_116_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_115_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_114_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_113_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_112_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_111_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_110_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_109_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_108_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_107_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_106_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_105_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_104_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_103_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_102_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_101_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_100_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_99_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_98_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_97_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_96_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_95_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_94_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_93_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_92_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_91_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_90_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_89_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_88_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_87_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_86_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_85_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_84_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_83_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_82_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_81_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_80_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_79_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_78_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_77_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_76_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_75_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_74_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_73_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_72_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_71_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_70_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_69_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_68_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_67_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_66_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_65_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_64_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_63_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_62_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_61_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_60_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_59_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_58_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_57_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_56_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_55_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_54_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_53_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_52_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_51_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_50_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_49_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_48_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_47_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_46_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_45_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_44_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_43_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_42_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_41_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_40_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_39_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_38_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_37_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_36_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_35_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_34_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_33_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_32_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_31_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_30_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_29_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_28_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_27_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_26_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_25_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_24_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_23_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_22_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_21_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_20_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_19_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_18_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_17_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_16_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_15_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_14_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_13_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_12_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_11_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_10_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_9_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_8_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_7_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_6_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_5_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_4_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_3_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_2_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_1_N3,
         Inst_forkAE_CipherInst_RF_RS2_SFF_0_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_127_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_126_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_125_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_124_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_123_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_122_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_121_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_120_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_119_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_118_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_117_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_116_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_115_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_114_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_113_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_112_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_111_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_110_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_109_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_108_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_107_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_106_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_105_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_104_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_103_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_102_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_101_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_100_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_99_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_98_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_97_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_96_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_95_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_94_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_93_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_92_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_91_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_90_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_89_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_88_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_87_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_86_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_85_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_84_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_83_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_82_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_81_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_80_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_79_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_78_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_77_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_76_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_75_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_74_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_73_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_72_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_71_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_70_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_69_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_68_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_67_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_66_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_65_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_64_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_63_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_62_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_61_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_60_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_59_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_58_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_57_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_56_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_55_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_54_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_53_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_52_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_51_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_50_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_49_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_48_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_47_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_46_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_45_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_44_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_43_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_42_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_41_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_40_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_39_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_38_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_37_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_36_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_35_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_34_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_33_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_32_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_31_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_30_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_29_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_28_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_27_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_26_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_25_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_24_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_23_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_22_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_21_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_20_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_19_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_18_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_17_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_16_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_15_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_14_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_13_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_12_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_11_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_10_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_9_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_8_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_7_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_6_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_5_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_4_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_3_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_2_N3,
         Inst_forkAE_CipherInst_RF_RS1_SFF_1_N3, n1, n2, n3, n4, n5, n6, n7,
         n8, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5718, n5719, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213;
  wire   [5:2] Inst_forkAE_CipherInst_ROUND_CST;
  wire   [127:0] Inst_forkAE_MainPart1_Auth_Reg_Output;
  wire   [127:0] Inst_forkAE_MainPart2_Auth_Reg_Output;
  wire   [127:0] Inst_forkAE_CipherInst_RF_S_MID_D2;
  wire   [127:0] Inst_forkAE_CipherInst_RF_S_MID_D1;
  wire   [63:2] Inst_forkAE_CipherInst_RF_SHIFT2_OUT;
  wire   [15:10] Inst_forkAE_CipherInst_RF_SHIFT1_OUT;
  wire   [124:8] Inst_forkAE_CipherInst_RF_S_MID_C1;
  wire   [124:64] Inst_forkAE_CipherInst_RF_S_MID_C2;
  wire   [127:0] Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv;

  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_23_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_62_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(n3), .QN(n484) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_2_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_49_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .QN(n465) );
  SEDFFTRX2 Inst_forkAE_CipherInst_CL_STATE_reg_2_ ( .RN(
        Inst_forkAE_ControlInst_fsm_state_1_), .D(
        Inst_forkAE_CipherInst_ROUND_CST[2]), .E(Inst_forkAE_CipherInst_LAST), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .QN(Inst_forkAE_CipherInst_CL_n27) );
  SEDFFTRX2 Inst_forkAE_CipherInst_CL_STATE_reg_4_ ( .RN(
        Inst_forkAE_ControlInst_fsm_state_1_), .D(
        Inst_forkAE_CipherInst_ROUND_CST[4]), .E(Inst_forkAE_CipherInst_LAST), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n6), .QN(
        Inst_forkAE_CipherInst_CL_n23) );
  SEDFFTRX2 Inst_forkAE_CipherInst_CL_STATE_reg_5_ ( .RN(
        Inst_forkAE_ControlInst_fsm_state_1_), .D(
        Inst_forkAE_CipherInst_ROUND_CST[5]), .E(Inst_forkAE_CipherInst_LAST), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n4), .QN(
        Inst_forkAE_CipherInst_CL_n22) );
  TLATNX2 Inst_forkAE_CipherInst_KE_CLK_GATE_K_reg ( .D(
        Inst_forkAE_CipherInst_KE_N2), .GN(clk), .QN(n462) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_22_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_61_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_62_), .QN(n483) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_21_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_60_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_61_), .QN(n482) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_20_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_59_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_60_), .QN(n481) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_19_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_58_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_59_), .QN(n480) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_18_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_57_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_58_), .QN(n479) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_17_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_56_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_57_), .QN(n478) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_16_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_7_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_56_), .QN(n477) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_15_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_6_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_7_), .QN(n476) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_14_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_5_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_6_), .QN(n475) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_13_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_4_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_5_), .QN(n474) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_12_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_3_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_4_), .QN(n473) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_11_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_2_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_3_), .QN(n472) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_10_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_1_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_2_), .QN(n471) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_9_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_0_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_1_), .QN(n470) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_8_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_55_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_0_), .QN(n469) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_7_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_54_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_55_), .QN(n468) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_6_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_53_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_54_), .QN(n467) );
  SEDFFTRX2 Inst_forkAE_LFSRInst_Reg_reg_5_ ( .RN(n5715), .D(
        Inst_forkAE_CipherInst_TK1_DEC_52_), .E(done), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .Q(Inst_forkAE_CipherInst_TK1_DEC_53_), .QN(n466) );
  SDFFTRXL Inst_forkAE_CipherInst_CL_COUNTER_reg_1_ ( .RN(
        Inst_forkAE_CipherInst_CL_n34), .D(n5719), .SI(1'b0), .SE(1'b0), .CK(
        clk), .Q(n2), .QN(n463) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_96_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_96_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_16_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_32_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_32_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_96_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_14_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_14_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_78_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_1_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_1_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_65_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_124_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_124_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_52_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_120_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_120_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_48_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_116_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_116_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_4_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_112_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_112_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_0_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_108_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_108_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_60_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_104_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_104_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_56_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_100_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_100_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_20_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_92_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_92_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_44_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_84_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_84_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_12_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_76_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_76_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_28_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_68_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_68_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_36_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_62_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_62_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_126_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_61_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_61_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_125_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_60_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_60_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_124_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_59_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_59_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_123_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_58_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_58_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_122_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_57_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_57_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_121_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_56_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_56_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_120_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_54_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_54_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_118_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_53_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_53_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_117_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_52_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_52_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_116_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_51_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_51_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_115_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_50_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_50_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_114_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_49_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_49_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_113_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_48_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_48_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_112_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_46_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_46_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_110_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_45_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_45_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_109_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_44_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_44_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_108_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_43_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_43_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_107_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_42_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_42_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_106_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_41_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_41_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_105_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_40_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_40_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_104_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_38_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_38_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_102_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_37_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_37_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_101_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_36_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_36_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_100_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_35_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_35_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_99_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_34_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_34_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_98_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_33_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_33_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_97_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_30_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_30_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_94_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_29_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_29_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_93_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_28_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_28_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_92_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_27_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_27_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_91_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_26_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_26_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_90_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_25_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_25_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_89_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_24_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_24_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_88_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_22_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_22_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_86_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_21_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_21_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_85_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_20_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_20_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_84_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_19_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_19_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_83_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_18_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_18_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_82_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_17_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_17_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_81_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_16_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_16_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_80_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_13_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_13_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_77_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_12_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_12_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_76_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_11_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_11_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_75_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_10_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_10_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_74_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_9_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_9_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_73_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_8_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_8_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_72_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_6_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_6_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_70_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_5_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_5_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_69_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_4_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_4_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_68_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_3_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_3_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_67_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_2_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_2_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_66_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_0_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_0_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_64_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_124_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_124_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_52_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_116_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_116_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_4_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_112_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_112_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_0_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_108_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_108_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_60_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_104_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_104_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_56_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_62_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_62_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_126_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_61_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_61_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_125_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_60_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_60_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_124_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_59_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_59_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_123_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_58_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_58_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_122_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_57_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_57_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_121_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_56_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_56_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_120_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_54_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_54_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_118_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_53_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_53_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_117_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_52_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_52_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_116_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_51_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_51_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_115_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_50_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_50_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_114_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_49_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_49_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_113_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_48_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_48_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_112_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_46_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_46_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_110_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_45_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_45_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_109_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_44_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_44_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_108_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_43_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_43_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_107_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_42_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_42_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_106_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_41_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_41_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_105_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_40_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_40_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_104_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_38_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_38_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_102_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_37_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_37_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_101_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_36_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_36_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_100_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_35_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_35_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_99_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_34_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_34_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_98_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_33_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_33_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_97_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_32_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_32_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_96_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_30_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_30_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_94_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_29_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_29_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_93_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_28_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_28_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_92_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_27_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_27_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_91_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_26_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_26_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_90_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_25_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_25_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_89_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_24_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_24_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_88_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_22_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_22_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_86_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_21_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_21_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_85_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_20_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_20_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_84_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_19_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_19_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_83_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_18_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_18_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_82_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_17_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_17_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_81_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_16_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_16_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_80_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_14_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_14_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_78_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_13_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_13_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_77_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_12_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_12_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_76_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_11_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_11_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_75_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_10_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_10_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_74_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_9_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_9_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_73_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_8_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_8_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_72_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_6_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_6_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_70_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_5_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_5_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_69_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_4_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_4_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_68_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_3_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_3_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_67_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_2_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_2_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_66_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_1_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_1_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_65_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_0_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_0_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_64_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_112_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_112_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[0]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_104_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_104_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[56]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_82_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_82_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[10]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_16_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_16_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[80]) );
  SEDFFTRX2 Inst_forkAE_CipherInst_CL_STATE_reg_1_ ( .RN(
        Inst_forkAE_ControlInst_fsm_state_1_), .D(n5718), .E(
        Inst_forkAE_CipherInst_LAST), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n464)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_36_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_36_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[100]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_62_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_62_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[126]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_61_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_61_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[125]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_60_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_60_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[124]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_59_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_59_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[123]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_58_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_58_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[122]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_57_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_57_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[121]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_56_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_56_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[120]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_55_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_55_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[119]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_54_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_54_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[118]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_53_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_53_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[117]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_52_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_52_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[116]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_50_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_50_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[114]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_49_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_49_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[113]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_7_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_7_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[71]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_6_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_6_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[70]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_5_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_5_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[69]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_4_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_4_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[68]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_3_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_3_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[67]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_2_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_2_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[66]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_1_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_1_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[65]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_0_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_0_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[64]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_48_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_48_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[112]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_42_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_42_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[106]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_40_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_40_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[104]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_34_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_34_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[98]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_33_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_33_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[97]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_26_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_26_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[90]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_25_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_25_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[89]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_15_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_15_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[79]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_14_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_14_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[78]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_13_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_13_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[77]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_11_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_11_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[75]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_63_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_63_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[127]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_51_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_51_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[115]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_47_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_47_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[111]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_46_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_46_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[110]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_45_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_45_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[109]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_44_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_44_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[108]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_43_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_43_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[107]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_41_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_41_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[105]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_32_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_32_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_31_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_31_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[95]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_30_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_30_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[94]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_29_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_29_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[93]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_28_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_28_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[92]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_27_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_27_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[91]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_24_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_24_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[88]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_12_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_12_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[76]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_9_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_9_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[73]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_39_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_39_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[103]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_38_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_38_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[102]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_37_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_37_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[101]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_35_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_35_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[99]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_23_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_23_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[87]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_22_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_22_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[86]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_21_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_21_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[85]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_19_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_19_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[83]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_20_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_20_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[84]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_10_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_10_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[74]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_8_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_8_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[72]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_124_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_124_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[52]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_116_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_116_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[4]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_108_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_108_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[60]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_13_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n273), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[13]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_17_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n277), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[17]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_21_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n281), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[21]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_32_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n292), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[32]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_36_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n296), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[36]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_40_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n300), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[40]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_44_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n304), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[44]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_48_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n308), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[48]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_52_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n312), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[52]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_56_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n316), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[56]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_60_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n320), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[60]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_65_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n325), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[65]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_73_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n333), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[73]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_81_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n341), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[81]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_89_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n349), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[89]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_96_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n356), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[96]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_100_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n360), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[100]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_104_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n364), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[104]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_108_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n368), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[108]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_112_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n372), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[112]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_116_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n376), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[116]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_120_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n380), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[120]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_124_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n384), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[124]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_66_ ( .D(n7768), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[66]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_69_ ( .D(n7771), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[69]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_74_ ( .D(n7776), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[74]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_77_ ( .D(n7779), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[77]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_82_ ( .D(n7784), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[82]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_85_ ( .D(n7787), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[85]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_87_ ( .D(n7789), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[87]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_90_ ( .D(n7792), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[90]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_93_ ( .D(n7795), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[93]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_95_ ( .D(n7797), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[95]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_96_ ( .D(n7798), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_17_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_17_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[81]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_18_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_18_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[82]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_1_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n261), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[1]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_6_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n266), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[6]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_14_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n274), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[14]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_22_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n282), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[22]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_30_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n290), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[30]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_33_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n293), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[33]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_37_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n297), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[37]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_38_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n298), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[38]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_41_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n301), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[41]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_45_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n305), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[45]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_46_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n306), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[46]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_49_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n309), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[49]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_53_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n313), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[53]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_54_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n314), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[54]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_57_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n317), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[57]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_61_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n321), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[61]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_62_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n322), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[62]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_70_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n330), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[70]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_78_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n338), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[78]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_86_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n346), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[86]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_94_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n354), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[94]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_97_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n357), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[97]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_101_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n361), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[101]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_102_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n362), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[102]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_105_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n365), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[105]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_109_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n369), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[109]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_110_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n370), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[110]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_113_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n373), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[113]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_117_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n377), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[117]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_118_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n378), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[118]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_121_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n381), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[121]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_125_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n385), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[125]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_126_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n386), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[126]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_1_ ( .D(n7703), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[1]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_6_ ( .D(n7708), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[6]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_9_ ( .D(n7711), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[9]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_14_ ( .D(n7716), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[14]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_22_ ( .D(n7724), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[22]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_25_ ( .D(n7727), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[25]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_30_ ( .D(n7732), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[30]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_33_ ( .D(n7735), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[33]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_37_ ( .D(n7739), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[37]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_38_ ( .D(n7740), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[38]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_41_ ( .D(n7743), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[41]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_45_ ( .D(n7747), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[45]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_46_ ( .D(n7748), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[46]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_49_ ( .D(n7751), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[49]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_53_ ( .D(n7755), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[53]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_54_ ( .D(n7756), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[54]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_57_ ( .D(n7759), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[57]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_61_ ( .D(n7763), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[61]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_62_ ( .D(n7764), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[62]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_97_ ( .D(n7799), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[97]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_101_ ( .D(n7803), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[101]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_102_ ( .D(n7804), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[102]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_105_ ( .D(n7807), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[105]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_109_ ( .D(n7811), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[109]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_110_ ( .D(n7812), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[110]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_113_ ( .D(n7815), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[113]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_117_ ( .D(n7819), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[117]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_118_ ( .D(n7820), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[118]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_121_ ( .D(n7823), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[121]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_125_ ( .D(n7827), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[125]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_126_ ( .D(n7828), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[126]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_82_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_82_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_10_) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_127_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n387), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[127]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_127_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_127_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_55_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_125_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_125_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_53_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_123_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_123_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_51_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_122_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_122_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_50_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_119_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_119_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_7_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_117_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_117_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_5_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_115_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_115_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_3_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_114_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_114_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_2_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_111_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_111_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_63_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_109_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_109_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_61_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_107_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_107_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_59_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_106_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_106_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_58_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_101_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_101_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_21_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_98_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_98_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_18_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_93_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_93_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_45_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_90_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_90_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_42_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_89_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_89_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_41_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_85_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_85_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_13_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_82_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_82_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_10_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_81_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_81_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_9_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_77_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_77_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_29_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_74_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_74_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_26_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_73_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_73_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_25_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_69_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_69_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_37_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_66_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_66_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_34_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_63_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_63_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_127_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_55_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_55_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_119_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_47_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_47_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_111_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_39_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_39_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_103_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_31_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_31_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_95_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_15_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_15_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_79_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_7_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_7_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_71_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_127_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_127_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_55_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_125_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_125_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_53_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_123_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_123_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_51_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_122_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_122_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_50_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_121_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_121_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_49_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_120_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_120_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_48_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_119_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_119_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_7_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_117_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_117_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_5_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_115_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_115_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_3_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_114_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_114_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_2_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_113_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_113_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_1_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_111_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_111_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_63_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_109_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_109_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_61_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_107_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_107_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_59_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_106_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_106_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_58_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_105_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_105_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_57_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_103_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_103_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_23_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_101_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_101_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_21_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_100_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_100_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_20_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_99_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_99_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_19_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_98_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_98_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_18_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_97_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_97_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_17_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_96_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_96_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_16_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_95_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_95_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_47_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_93_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_93_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_45_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_92_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_92_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_44_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_91_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_91_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_43_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_90_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_90_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_42_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_89_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_89_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_41_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_88_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_88_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_40_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_87_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_87_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_15_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_85_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_85_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_13_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_84_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_84_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_12_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_83_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_83_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_11_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_81_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_81_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_9_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_80_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_80_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_8_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_79_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_79_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_31_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_77_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_77_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_29_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_76_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_76_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_28_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_75_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_75_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_27_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_74_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_74_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_26_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_73_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_73_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_25_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_72_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_72_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_24_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_71_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_71_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_39_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_69_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_69_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_37_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_68_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_68_N3), .SI(1'b0), .SE(1'b0), .CK(
        n428), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_36_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_67_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_67_N3), .SI(1'b0), .SE(1'b0), .CK(
        n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_35_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_66_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_66_N3), .SI(1'b0), .SE(1'b0), .CK(
        n430), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_34_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_65_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_65_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_33_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_64_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_64_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_32_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_63_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_63_N3), .SI(1'b0), .SE(1'b0), .CK(
        n434), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_127_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_55_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_55_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_119_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_47_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_47_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_111_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_39_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_39_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_103_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_31_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_31_N3), .SI(1'b0), .SE(1'b0), .CK(
        n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_95_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_23_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_23_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_87_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_15_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_15_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_79_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_7_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_7_N3), .SI(1'b0), .SE(1'b0), .CK(
        n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_71_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_65_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_65_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_33_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_23_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_23_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_87_) );
  SDFFSQXL Inst_forkAE_LFSRInst_Reg_reg_3_ ( .D(Inst_forkAE_LFSRInst_n62), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CipherInst_TK1_DEC_51_) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_2_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n262), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[2]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_3_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n263), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[3]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_5_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n265), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[5]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_7_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n267), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[7]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_10_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n270), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[10]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_11_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n271), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[11]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_15_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n275), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[15]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_18_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n278), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[18]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_19_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n279), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[19]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_23_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n283), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[23]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_26_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n286), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[26]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_27_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n287), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[27]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_29_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n289), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[29]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_31_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n291), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[31]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_34_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n294), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[34]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_35_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n295), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[35]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_39_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n299), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[39]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_42_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n302), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[42]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_43_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n303), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[43]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_47_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n307), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[47]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_50_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n310), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[50]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_51_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n311), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[51]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_55_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n315), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[55]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_58_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n318), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[58]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_59_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n319), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[59]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_63_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n323), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[63]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_66_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n326), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[66]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_67_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n327), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[67]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_69_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n329), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[69]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_71_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n331), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[71]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_74_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n334), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[74]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_75_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n335), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[75]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_77_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n337), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[77]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_79_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n339), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[79]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_82_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n342), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[82]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_83_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n343), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[83]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_85_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n345), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[85]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_87_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n347), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[87]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_90_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n350), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[90]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_91_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n351), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[91]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_93_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n353), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[93]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_95_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n355), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[95]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_98_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n358), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[98]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_99_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n359), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[99]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_103_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n363), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[103]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_106_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n366), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[106]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_107_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n367), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[107]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_111_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n371), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[111]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_114_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n374), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[114]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_115_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n375), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[115]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_119_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n379), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[119]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_122_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n382), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[122]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_123_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n383), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[123]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_2_ ( .D(n7704), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[2]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_3_ ( .D(n7705), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[3]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_5_ ( .D(n7707), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[5]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_7_ ( .D(n7709), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[7]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_10_ ( .D(n7712), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[10]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_11_ ( .D(n7713), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[11]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_13_ ( .D(n7715), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[13]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_15_ ( .D(n7717), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[15]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_17_ ( .D(n7719), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[17]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_18_ ( .D(n7720), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[18]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_19_ ( .D(n7721), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[19]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_21_ ( .D(n7723), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[21]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_23_ ( .D(n7725), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[23]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_26_ ( .D(n7728), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[26]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_27_ ( .D(n7729), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[27]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_29_ ( .D(n7731), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[29]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_31_ ( .D(n7733), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[31]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_32_ ( .D(n7734), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[32]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_34_ ( .D(n7736), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[34]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_35_ ( .D(n7737), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[35]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_36_ ( .D(n7738), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[36]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_39_ ( .D(n7741), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[39]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_40_ ( .D(n7742), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[40]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_42_ ( .D(n7744), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[42]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_43_ ( .D(n7745), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[43]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_44_ ( .D(n7746), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[44]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_47_ ( .D(n7749), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[47]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_48_ ( .D(n7750), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[48]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_50_ ( .D(n7752), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[50]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_51_ ( .D(n7753), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[51]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_52_ ( .D(n7754), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[52]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_55_ ( .D(n7757), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[55]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_56_ ( .D(n7758), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[56]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_58_ ( .D(n7760), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[58]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_59_ ( .D(n7761), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[59]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_60_ ( .D(n7762), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[60]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_63_ ( .D(n7765), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[63]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_65_ ( .D(n7767), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[65]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_67_ ( .D(n7769), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[67]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_71_ ( .D(n7773), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[71]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_73_ ( .D(n7775), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[73]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_75_ ( .D(n7777), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[75]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_79_ ( .D(n7781), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[79]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_81_ ( .D(n7783), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[81]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_83_ ( .D(n7785), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[83]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_89_ ( .D(n7791), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[89]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_91_ ( .D(n7793), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[91]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_98_ ( .D(n7800), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[98]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_99_ ( .D(n7801), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[99]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_100_ ( .D(n7802), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[100]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_103_ ( .D(n7805), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[103]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_104_ ( .D(n7806), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[104]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_106_ ( .D(n7808), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[106]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_107_ ( .D(n7809), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[107]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_108_ ( .D(n7810), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[108]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_111_ ( .D(n7813), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[111]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_112_ ( .D(n7814), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[112]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_114_ ( .D(n7816), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[114]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_115_ ( .D(n7817), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[115]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_116_ ( .D(n7818), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[116]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_119_ ( .D(n7821), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[119]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_120_ ( .D(n7822), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[120]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_122_ ( .D(n7824), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[122]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_123_ ( .D(n7825), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[123]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_124_ ( .D(n7826), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[124]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_127_ ( .D(n7829), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[127]) );
  SDFFSQXL Inst_forkAE_ControlInst_encdec_started_reg ( .D(
        Inst_forkAE_ControlInst_n31), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_ControlInst_encdec_started) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_0_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n260), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[0]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_4_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n264), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[4]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_8_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n268), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[8]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_9_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n269), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[9]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_12_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n272), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[12]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_16_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n276), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[16]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_20_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n280), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[20]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_24_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n284), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[24]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_25_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n285), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[25]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_28_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n288), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[28]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_64_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n324), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[64]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_68_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n328), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[68]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_72_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n332), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[72]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_76_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n336), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[76]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_80_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n340), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[80]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_84_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n344), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[84]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_88_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n348), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[88]) );
  SDFFSQXL Inst_forkAE_MainPart1_AuthRegInst_Output_reg_92_ ( .D(
        Inst_forkAE_MainPart1_AuthRegInst_n352), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_MainPart1_Auth_Reg_Output[92]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_0_ ( .D(n7702), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[0]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_4_ ( .D(n7706), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[4]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_8_ ( .D(n7710), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[8]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_12_ ( .D(n7714), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[12]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_16_ ( .D(n7718), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[16]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_20_ ( .D(n7722), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[20]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_24_ ( .D(n7726), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[24]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_28_ ( .D(n7730), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[28]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_64_ ( .D(n7766), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[64]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_68_ ( .D(n7770), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[68]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_70_ ( .D(n7772), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[70]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_72_ ( .D(n7774), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[72]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_76_ ( .D(n7778), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[76]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_78_ ( .D(n7780), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[78]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_80_ ( .D(n7782), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[80]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_84_ ( .D(n7786), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[84]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_86_ ( .D(n7788), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[86]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_88_ ( .D(n7790), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[88]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_92_ ( .D(n7794), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[92]) );
  SDFFSQXL Inst_forkAE_MainPart2_AuthRegInst_Output_reg_94_ ( .D(n7796), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Auth_Reg_Output[94]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_88_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_88_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_40_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_72_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_72_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_24_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_64_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_64_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_32_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_106_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_106_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[58]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_98_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_98_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[18]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_97_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_97_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[17]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_89_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_89_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[41]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_84_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_84_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[12]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_81_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_81_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[9]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_79_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_79_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[31]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_78_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_78_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[30]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_77_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_77_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[29]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_75_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_75_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[27]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_72_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_72_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[24]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_125_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_125_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[120]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_117_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_117_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[112]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_8_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N11), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_8_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_10_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N13), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_10_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_12_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N15), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_12_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_14_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N17), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_14_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_8_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N11), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_8_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_9_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N12), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_9_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_10_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N13), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_10_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_11_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N14), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_11_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_12_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N15), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_12_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_14_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N17), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_14_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_27_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N30), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_27_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_29_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N32), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_29_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_31_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N34), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_31_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_2_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N5), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_2_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_24_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N27), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_24_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_1_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N4), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_1_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_2_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N5), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_2_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_4_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N7), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_4_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_5_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N8), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_5_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_7_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N10), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_7_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_13_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N16), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_13_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_15_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N18), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_15_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_16_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N19), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_16_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_17_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N20), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_17_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_18_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N21), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_18_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_19_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N22), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_19_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_20_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N23), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_20_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_21_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N24), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_21_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_22_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N25), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_22_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_23_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N26), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_23_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_24_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N27), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_24_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_25_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N28), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_25_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_26_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N29), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_26_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_28_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N31), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_28_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_30_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N33), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_30_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_0_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N3), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_0_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_1_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N4), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_1_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_3_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N6), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_3_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_4_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N7), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_4_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_5_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N8), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_5_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_6_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N9), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_6_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_7_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N10), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_7_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_9_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N12), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_9_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_11_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N14), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_11_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_13_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N16), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_13_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_15_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N18), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_15_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_16_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N19), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_16_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_17_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N20), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_17_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_18_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N21), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_18_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_19_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N22), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_19_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_20_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N23), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_20_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_21_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N24), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_21_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_22_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N25), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_22_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_23_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N26), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_23_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_25_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N28), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_25_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_26_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N29), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_26_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_27_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N30), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_27_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_28_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N31), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_28_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_29_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N32), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_29_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_30_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N33), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_30_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX1_Output_reg_31_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX1_N34), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX1_31_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_0_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N3), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_0_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_3_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N6), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_3_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS_EX2_Output_reg_6_ ( .D(
        Inst_forkAE_CipherInst_RF_RS_EX2_N9), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_STATE_EX2_6_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_90_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_90_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[42]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_103_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_103_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[23]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_102_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_102_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[22]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_101_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_101_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[21]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_99_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_99_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[19]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_96_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_96_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[16]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_120_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_120_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[48]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_88_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_88_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[40]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_74_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_74_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[26]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_73_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_73_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[25]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_66_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_66_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[34]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_65_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_65_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[33]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_100_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_100_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[20]) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_0_ ( .D(n8086), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_0_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_1_ ( .D(n8087), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_1_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_2_ ( .D(n8088), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_2_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_3_ ( .D(n8089), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_3_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_4_ ( .D(n8090), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_4_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_5_ ( .D(n8091), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_5_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_6_ ( .D(n8092), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_6_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_8_ ( .D(n8094), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_8_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_9_ ( .D(n8095), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_9_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_10_ ( .D(n8096), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_10_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_11_ ( .D(n8097), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_11_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_12_ ( .D(n8098), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_12_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_13_ ( .D(n8099), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_13_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_14_ ( .D(n8100), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_14_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_16_ ( .D(n8102), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_16_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_17_ ( .D(n8103), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_17_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_18_ ( .D(n8104), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_18_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_19_ ( .D(n8105), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_19_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_20_ ( .D(n8106), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_20_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_21_ ( .D(n8107), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_21_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_22_ ( .D(n8108), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_22_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_24_ ( .D(n8110), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_24_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_25_ ( .D(n8111), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_25_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_26_ ( .D(n8112), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_26_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_27_ ( .D(n8113), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_27_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_28_ ( .D(n8114), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_28_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_29_ ( .D(n8115), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_29_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_30_ ( .D(n8116), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_30_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_32_ ( .D(n8118), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_32_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_33_ ( .D(n8119), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_33_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_34_ ( .D(n8120), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_34_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_35_ ( .D(n8121), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_35_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_36_ ( .D(n8122), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_36_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_37_ ( .D(n8123), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_37_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_38_ ( .D(n8124), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_38_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_40_ ( .D(n8126), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_40_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_41_ ( .D(n8127), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_41_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_42_ ( .D(n8128), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_42_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_43_ ( .D(n8129), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_43_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_44_ ( .D(n8130), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_44_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_45_ ( .D(n8131), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_45_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_46_ ( .D(n8132), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_46_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_48_ ( .D(n8134), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_48_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_49_ ( .D(n8135), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_49_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_50_ ( .D(n8136), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_50_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_51_ ( .D(n8137), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_51_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_52_ ( .D(n8138), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_52_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_53_ ( .D(n8139), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_53_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_54_ ( .D(n8140), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_54_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_56_ ( .D(n8142), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_56_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_57_ ( .D(n8143), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_57_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_58_ ( .D(n8144), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_58_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_59_ ( .D(n8145), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_59_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_60_ ( .D(n8146), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_60_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_61_ ( .D(n8147), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_61_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_62_ ( .D(n8148), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_62_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_64_ ( .D(n8150), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_64_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_65_ ( .D(n8151), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_65_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_66_ ( .D(n8152), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_66_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_67_ ( .D(n8153), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_67_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_68_ ( .D(n8154), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_68_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_69_ ( .D(n8155), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_69_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_70_ ( .D(n8156), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_70_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_72_ ( .D(n8158), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_72_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_73_ ( .D(n8159), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_73_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_74_ ( .D(n8160), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_74_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_75_ ( .D(n8161), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_75_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_76_ ( .D(n8162), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_76_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_77_ ( .D(n8163), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_77_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_78_ ( .D(n8164), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_78_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_80_ ( .D(n8166), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_80_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_81_ ( .D(n8167), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_81_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_82_ ( .D(n8168), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_82_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_83_ ( .D(n8169), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_83_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_84_ ( .D(n8170), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_84_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_85_ ( .D(n8171), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_85_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_86_ ( .D(n8172), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_86_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_88_ ( .D(n8174), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_88_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_89_ ( .D(n8175), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_89_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_90_ ( .D(n8176), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_90_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_91_ ( .D(n8177), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_91_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_92_ ( .D(n8178), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_92_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_93_ ( .D(n8179), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_93_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_94_ ( .D(n8180), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_94_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_96_ ( .D(n8182), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_96_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_97_ ( .D(n8183), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_97_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_98_ ( .D(n8184), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_98_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_99_ ( .D(n8185), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_99_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_100_ ( .D(n8186), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_100_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_101_ ( .D(n8187), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_101_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_102_ ( .D(n8188), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_102_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_104_ ( .D(n8190), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_104_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_105_ ( .D(n8191), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_105_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_106_ ( .D(n8192), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_106_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_107_ ( .D(n8193), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_107_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_108_ ( .D(n8194), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_108_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_109_ ( .D(n8195), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_109_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_110_ ( .D(n8196), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_110_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_112_ ( .D(n8198), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_112_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_113_ ( .D(n8199), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_113_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_114_ ( .D(n8200), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_114_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_115_ ( .D(n8201), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_115_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_116_ ( .D(n8202), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_116_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_117_ ( .D(n8203), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_117_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_118_ ( .D(n8204), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_118_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_120_ ( .D(n8206), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_120_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_121_ ( .D(n8207), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_121_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_122_ ( .D(n8208), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_122_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_123_ ( .D(n8209), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_123_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_124_ ( .D(n8210), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_124_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_125_ ( .D(n8211), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_125_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_126_ ( .D(n8212), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_126_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_0_ ( .D(n7318), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_0_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_1_ ( .D(n7319), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_1_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_2_ ( .D(n7320), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_2_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_3_ ( .D(n7321), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_3_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_4_ ( .D(n7322), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_4_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_5_ ( .D(n7323), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_5_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_6_ ( .D(n7324), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_6_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_8_ ( .D(n7326), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_8_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_9_ ( .D(n7327), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_9_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_10_ ( .D(n7328), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_10_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_11_ ( .D(n7329), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_11_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_12_ ( .D(n7330), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_12_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_13_ ( .D(n7331), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_13_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_14_ ( .D(n7332), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_14_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_16_ ( .D(n7334), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_16_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_17_ ( .D(n7335), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_17_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_18_ ( .D(n7336), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_18_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_19_ ( .D(n7337), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_19_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_20_ ( .D(n7338), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_20_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_21_ ( .D(n7339), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_21_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_22_ ( .D(n7340), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_22_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_24_ ( .D(n7342), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_24_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_25_ ( .D(n7343), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_25_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_26_ ( .D(n7344), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_26_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_27_ ( .D(n7345), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_27_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_28_ ( .D(n7346), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_28_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_29_ ( .D(n7347), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_29_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_30_ ( .D(n7348), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_30_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_32_ ( .D(n7350), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_32_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_33_ ( .D(n7351), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_33_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_34_ ( .D(n7352), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_34_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_35_ ( .D(n7353), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_35_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_36_ ( .D(n7354), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_36_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_37_ ( .D(n7355), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_37_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_38_ ( .D(n7356), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_38_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_40_ ( .D(n7358), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_40_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_41_ ( .D(n7359), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_41_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_42_ ( .D(n7360), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_42_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_43_ ( .D(n7361), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_43_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_44_ ( .D(n7362), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_44_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_45_ ( .D(n7363), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_45_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_46_ ( .D(n7364), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_46_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_48_ ( .D(n7366), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_48_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_49_ ( .D(n7367), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_49_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_50_ ( .D(n7368), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_50_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_51_ ( .D(n7369), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_51_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_52_ ( .D(n7370), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_52_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_53_ ( .D(n7371), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_53_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_54_ ( .D(n7372), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_54_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_56_ ( .D(n7374), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_56_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_57_ ( .D(n7375), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_57_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_58_ ( .D(n7376), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_58_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_59_ ( .D(n7377), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_59_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_60_ ( .D(n7378), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_60_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_61_ ( .D(n7379), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_61_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_62_ ( .D(n7380), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_62_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_64_ ( .D(n7382), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_64_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_65_ ( .D(n7383), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_65_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_66_ ( .D(n7384), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_66_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_67_ ( .D(n7385), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_67_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_68_ ( .D(n7386), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_68_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_69_ ( .D(n7387), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_69_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_70_ ( .D(n7388), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_70_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_72_ ( .D(n7390), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_72_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_73_ ( .D(n7391), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_73_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_74_ ( .D(n7392), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_74_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_75_ ( .D(n7393), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_75_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_76_ ( .D(n7394), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_76_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_77_ ( .D(n7395), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_77_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_78_ ( .D(n7396), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_78_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_80_ ( .D(n7398), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_80_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_81_ ( .D(n7399), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_81_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_82_ ( .D(n7400), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_82_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_83_ ( .D(n7401), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_83_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_84_ ( .D(n7402), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_84_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_85_ ( .D(n7403), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_85_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_86_ ( .D(n7404), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_86_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_88_ ( .D(n7406), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_88_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_89_ ( .D(n7407), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_89_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_90_ ( .D(n7408), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_90_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_91_ ( .D(n7409), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_91_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_92_ ( .D(n7410), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_92_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_93_ ( .D(n7411), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_93_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_94_ ( .D(n7412), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_94_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_96_ ( .D(n7414), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_96_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_97_ ( .D(n7415), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_97_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_98_ ( .D(n7416), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_98_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_99_ ( .D(n7417), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_99_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_100_ ( .D(n7418), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_100_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_101_ ( .D(n7419), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_101_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_102_ ( .D(n7420), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_102_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_104_ ( .D(n7422), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_104_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_105_ ( .D(n7423), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_105_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_106_ ( .D(n7424), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_106_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_107_ ( .D(n7425), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_107_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_108_ ( .D(n7426), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_108_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_109_ ( .D(n7427), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_109_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_110_ ( .D(n7428), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_110_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_112_ ( .D(n7430), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_112_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_113_ ( .D(n7431), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_113_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_114_ ( .D(n7432), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_114_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_115_ ( .D(n7433), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_115_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_116_ ( .D(n7434), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_116_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_117_ ( .D(n7435), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_117_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_118_ ( .D(n7436), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_118_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_120_ ( .D(n7438), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_120_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_121_ ( .D(n7439), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_121_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_122_ ( .D(n7440), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_122_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_123_ ( .D(n7441), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_123_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_124_ ( .D(n7442), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_124_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_125_ ( .D(n7443), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_125_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_126_ ( .D(n7444), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_126_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_87_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_87_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[15]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_86_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_86_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[14]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_85_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_85_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[13]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_83_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_83_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[11]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_80_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_80_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[8]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_122_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_122_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[122]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_114_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_114_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[114]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_106_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_106_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[106]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_127_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_127_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[55]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_126_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_126_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[54]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_125_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_125_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[53]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_123_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_123_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[51]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_122_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_122_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[50]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_121_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_121_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[49]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_119_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_119_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[7]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_118_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_118_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[6]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_117_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_117_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[5]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_115_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_115_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[3]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_114_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_114_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[2]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_113_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_113_N3), .SI(1'b0), .SE(1'b0), .CK(
        n424), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[1]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_111_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_111_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[63]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_110_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_110_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[62]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_109_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_109_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[61]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_107_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_107_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[59]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_105_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_105_N3), .SI(1'b0), .SE(1'b0), .CK(
        n423), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[57]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_95_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_95_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[47]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_94_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_94_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[46]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_93_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_93_N3), .SI(1'b0), .SE(1'b0), .CK(
        n418), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[45]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_92_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_92_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[44]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_91_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_91_N3), .SI(1'b0), .SE(1'b0), .CK(
        n426), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[43]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_76_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_76_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[28]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_71_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_71_N3), .SI(1'b0), .SE(1'b0), .CK(
        n421), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[39]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_70_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_70_N3), .SI(1'b0), .SE(1'b0), .CK(
        n420), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[38]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_69_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_69_N3), .SI(1'b0), .SE(1'b0), .CK(
        n419), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[37]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_68_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_68_N3), .SI(1'b0), .SE(1'b0), .CK(
        n417), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[36]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_67_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_67_N3), .SI(1'b0), .SE(1'b0), .CK(
        n425), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[35]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS1_SFF_64_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS1_SFF_64_N3), .SI(1'b0), .SE(1'b0), .CK(
        n422), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[32]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_0_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_0_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[0]) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_7_ ( .D(n8093), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_7_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_15_ ( .D(n8101), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_15_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_23_ ( .D(n8109), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_23_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_31_ ( .D(n8117), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_31_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_39_ ( .D(n8125), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_39_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_47_ ( .D(n8133), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_47_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_55_ ( .D(n8141), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_55_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_63_ ( .D(n8149), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_63_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_71_ ( .D(n8157), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_71_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_79_ ( .D(n8165), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_79_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_87_ ( .D(n8173), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_87_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_95_ ( .D(n8181), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_95_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_103_ ( .D(n8189), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_103_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_111_ ( .D(n8197), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_111_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_119_ ( .D(n8205), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_119_) );
  SDFFSQXL Inst_forkAE_MainPart2_TagRegInst_Output_reg_127_ ( .D(n8213), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart2_Tag_Reg_Output_127_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_7_ ( .D(n7325), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_7_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_15_ ( .D(n7333), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_15_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_23_ ( .D(n7341), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_23_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_31_ ( .D(n7349), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_31_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_39_ ( .D(n7357), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_39_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_47_ ( .D(n7365), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_47_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_55_ ( .D(n7373), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_55_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_63_ ( .D(n7381), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_63_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_71_ ( .D(n7389), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_71_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_79_ ( .D(n7397), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_79_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_87_ ( .D(n7405), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_87_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_95_ ( .D(n7413), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_95_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_103_ ( .D(n7421), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_103_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_111_ ( .D(n7429), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_111_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_119_ ( .D(n7437), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_119_) );
  SDFFSQXL Inst_forkAE_MainPart1_TagRegInst_Output_reg_127_ ( .D(n7445), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_MainPart1_Tag_Reg_Output_127_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_124_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_124_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[124]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_116_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_116_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[116]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_108_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_108_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[108]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_100_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_100_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[100]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_124_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_124_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[124]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_120_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_120_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[120]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_116_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_116_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[116]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_112_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_112_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[112]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_108_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_108_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[108]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_104_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_104_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[104]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_100_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_100_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[100]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_80_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_80_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[80]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_72_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_72_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[72]) );
  SDFFSQXL Inst_forkAE_ControlInst_fsm_state_reg_0_ ( .D(
        Inst_forkAE_ControlInst_n33), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_ControlInst_fsm_state_0_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_126_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_126_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_54_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_118_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_118_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_6_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_110_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_110_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_62_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_102_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_102_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_22_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_126_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_126_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_54_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_118_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_118_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n433), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_6_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_110_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_110_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n435), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_62_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_102_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_102_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n432), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_22_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_94_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_94_N3), .SI(1'b0), .SE(1'b0), .CK(
        n429), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_46_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_86_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_86_N3), .SI(1'b0), .SE(1'b0), .CK(
        n431), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_14_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_78_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_78_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_30_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_1_SFF_70_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_1_SFF_70_N3), .SI(1'b0), .SE(1'b0), .CK(
        n427), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_38_) );
  SDFFSQXL Inst_forkAE_CipherInst_CL_STATE_reg_0_ ( .D(
        Inst_forkAE_CipherInst_CL_n44), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_forkAE_CipherInst_CL_STATE_0_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_126_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_126_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[124]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_118_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_118_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[116]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_110_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_110_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[108]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_109_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_109_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[104]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_103_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_103_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_23_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_121_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_121_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_49_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_113_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_113_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_1_)
         );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_105_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_105_N3), .SI(1'b0), .SE(1'b0), 
        .CK(n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_57_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_99_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_99_N3), .SI(1'b0), .SE(1'b0), .CK(
        n438), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_19_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_97_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_97_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_17_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_95_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_95_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_47_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_91_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_91_N3), .SI(1'b0), .SE(1'b0), .CK(
        n443), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_43_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_86_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_86_N3), .SI(1'b0), .SE(1'b0), .CK(
        n441), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_14_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_83_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_83_N3), .SI(1'b0), .SE(1'b0), .CK(
        n444), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_11_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_80_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_80_N3), .SI(1'b0), .SE(1'b0), .CK(
        n439), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_8_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_79_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_79_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_31_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_75_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_75_N3), .SI(1'b0), .SE(1'b0), .CK(
        n437), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_27_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_71_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_71_N3), .SI(1'b0), .SE(1'b0), .CK(
        n442), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_39_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_67_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_67_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_35_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_87_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_87_N3), .SI(1'b0), .SE(1'b0), .CK(
        n446), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_15_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_72_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_72_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[72]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_46_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_46_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[58]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_38_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_38_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[50]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_37_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_37_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[55]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_13_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_13_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[8]) );
  SDFFSQXL Inst_forkAE_LFSRInst_Reg_reg_0_ ( .D(n5716), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_TK1_DEC_48_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_122_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_122_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[122]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_114_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_114_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[114]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_106_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_106_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[106]) );
  SDFFSQXL Inst_forkAE_CipherInst_CL_COUNTER_reg_2_ ( .D(
        Inst_forkAE_CipherInst_CL_N15), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_forkAE_CipherInst_CL_COUNTER_2_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_98_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_98_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[98]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_98_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_98_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[98]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_58_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_58_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[58]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_50_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_50_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[50]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_42_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_42_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[42]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_34_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_34_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[34]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_58_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_58_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[58]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_50_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_50_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[50]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_42_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_42_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[42]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_34_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_34_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[34]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_121_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_121_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[121]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_113_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_113_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[113]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_105_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_105_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[105]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_113_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_113_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[113]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_105_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_105_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[105]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_120_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_120_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[120]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_112_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_112_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[112]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_104_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_104_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[104]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_64_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_64_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[64]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_0_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_0_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[0]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_96_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_96_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_24_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_24_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[24]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_97_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_97_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[97]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_97_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_97_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[97]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_9_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_9_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[9]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_59_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_59_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[59]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_51_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_51_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[51]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_43_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_43_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[43]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_35_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_35_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[35]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_123_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_123_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[123]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_115_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_115_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[115]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_107_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_107_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[107]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_49_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_49_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[49]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_101_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_101_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_125_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_125_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[120]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_117_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_117_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[112]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_109_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_109_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[104]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_59_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_59_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[59]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_43_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_43_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[43]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_35_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_35_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[35]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_99_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_99_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[99]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_127_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_127_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[127]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_119_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_119_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[119]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_111_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_111_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[111]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_103_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_103_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[103]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_101_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_101_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_123_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_123_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[123]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_115_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_115_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[115]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_107_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_107_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[107]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_63_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_63_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[63]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_57_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_57_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[57]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_55_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_55_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[55]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_49_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_49_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[49]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_47_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_47_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[47]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_41_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_41_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[41]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_39_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_39_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[39]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_33_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_33_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[33]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_102_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_102_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[100]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_88_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_88_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[88]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_80_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_80_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[80]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_64_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_64_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[64]) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_94_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_94_N3), .SI(1'b0), .SE(1'b0), .CK(
        n440), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_78_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_78_N3), .SI(1'b0), .SE(1'b0), .CK(
        n445), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_) );
  SDFFSQXL Inst_forkAE_CipherInst_KE_RS2_2_SFF_70_Q_reg ( .D(
        Inst_forkAE_CipherInst_KE_RS2_2_SFF_70_N3), .SI(1'b0), .SE(1'b0), .CK(
        n436), .SN(1'b1), .Q(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_62_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_62_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[42]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_54_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_54_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[34]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_13_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_13_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[23]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_99_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_99_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[99]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_51_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_51_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[51]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_15_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_15_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[15]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_45_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_45_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[63]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_61_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_61_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[47]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_53_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_53_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[39]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_29_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_29_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[24]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_21_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_21_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[16]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_66_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_66_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[66]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_74_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_74_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[74]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_90_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_90_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[90]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_82_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_82_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[82]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_121_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_121_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[121]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_90_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_90_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[90]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_82_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_82_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[82]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_74_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_74_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[74]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_66_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_66_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[66]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_2_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_2_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[2]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_2_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_2_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[2]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_61_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_61_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[56]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_91_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_91_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[91]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_83_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_83_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[83]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_75_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_75_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[75]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_67_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_67_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[67]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_53_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_53_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[48]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_45_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_45_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[40]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_37_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_37_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[32]) );
  SDFFSQXL Inst_forkAE_CipherInst_CL_COUNTER_reg_0_ ( .D(
        Inst_forkAE_CipherInst_CL_N13), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(Inst_forkAE_CipherInst_CL_COUNTER_0_) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_18_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_18_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[18]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_10_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_10_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[10]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_10_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_10_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[10]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_96_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_96_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[96]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_8_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_8_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[8]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_26_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_26_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[26]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_26_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_26_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[26]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_18_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_18_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[18]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_28_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_28_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[28]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_24_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_24_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[24]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_20_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_20_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[20]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_16_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_16_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[16]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_12_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_12_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[12]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_4_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_4_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[4]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_28_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_28_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[28]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_20_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_20_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[20]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_16_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_16_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[16]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_12_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_12_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[12]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_4_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_4_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[4]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_1_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_1_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[1]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_27_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_27_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[27]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_19_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_19_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[19]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_11_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_11_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[11]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_92_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_92_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[92]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_88_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_88_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[88]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_84_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_84_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[84]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_76_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_76_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[76]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_68_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_68_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[68]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_29_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_29_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_21_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_21_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_93_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_93_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[88]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_85_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_85_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[80]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_77_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_77_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[72]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_69_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_69_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[64]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_5_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_5_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_93_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_93_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[88]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_85_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_85_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[80]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_69_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_69_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[64]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_5_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_5_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_91_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_91_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[91]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_83_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_83_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[83]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_75_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_75_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[75]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_67_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_67_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[67]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_25_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_25_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[25]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_17_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_17_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[17]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_11_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_11_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[11]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_3_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_3_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[3]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_57_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_57_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[57]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_41_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_41_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[41]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_33_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_33_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[33]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_77_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_77_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[72]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_19_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_19_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[19]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_7_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_7_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[7]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_30_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_30_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_22_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_22_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_14_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_14_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_6_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_6_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_3_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_3_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[3]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_65_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_65_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[65]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_31_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_31_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[31]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_23_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_23_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[23]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_94_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_94_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[92]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_86_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_86_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[84]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_78_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_78_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[76]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_70_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_70_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C2[68]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_27_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_27_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[27]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_73_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_73_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[73]) );
  SDFFSX2 Inst_forkAE_LFSRInst_Reg_reg_4_ ( .D(Inst_forkAE_LFSRInst_n61), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CipherInst_TK1_DEC_52_), .QN(Inst_forkAE_LFSRInst_n51) );
  SDFFSX2 Inst_forkAE_LFSRInst_Reg_reg_1_ ( .D(Inst_forkAE_LFSRInst_n63), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CipherInst_TK1_DEC_49_), .QN(Inst_forkAE_LFSRInst_n52) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_89_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_89_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[89]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_81_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_81_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[81]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_8_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_8_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[8]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_60_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_60_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[60]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_56_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_56_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[56]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_44_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_44_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[44]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_40_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_40_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[40]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_36_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_36_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[36]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_32_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_32_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[32]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_52_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_52_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[52]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_119_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_119_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[119]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_111_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_111_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[111]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_92_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_92_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[92]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_84_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_84_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[84]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_76_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_76_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[76]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_68_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_68_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[68]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_95_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_95_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[95]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_87_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_87_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[87]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_79_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_79_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[79]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_9_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_9_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[9]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_1_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_1_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[1]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_89_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_89_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[89]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_81_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_81_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[81]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_65_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_65_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[65]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_71_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_71_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[71]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_25_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_25_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[25]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_17_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_17_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[17]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_73_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_73_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[73]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_32_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_32_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[32]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_56_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_56_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[56]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_52_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_52_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[52]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS2_SFF_48_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS2_SFF_48_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D2[48]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_60_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_60_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[60]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_44_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_44_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[44]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_40_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_40_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[40]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_36_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_36_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[36]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_103_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_103_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[103]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_118_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_118_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[116]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_110_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_110_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[108]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_126_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_126_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[124]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_48_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_48_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[48]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_102_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_102_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[100]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_127_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_127_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[127]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_63_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_63_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[63]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_55_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_55_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[55]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_47_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_47_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[47]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_7_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_7_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[7]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_6_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_6_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_62_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_62_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[60]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_54_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_54_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[52]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_46_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_46_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[44]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_38_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_38_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[36]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_94_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_94_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[92]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_86_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_86_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[84]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_78_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_78_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[76]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_70_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_70_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[68]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_22_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_22_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[20]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_14_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_14_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[12]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_15_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_15_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[15]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_39_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_39_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[39]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_23_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_23_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[23]) );
  SDFFSX2 Inst_forkAE_CipherInst_CL_STATE_reg_3_ ( .D(
        Inst_forkAE_CipherInst_CL_n43), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        1'b1), .Q(n461) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_95_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_95_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[95]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_87_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_87_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[87]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_79_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_79_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[79]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_31_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_31_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[31]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_30_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_30_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_C1[28]) );
  SDFFSQXL Inst_forkAE_CipherInst_RF_RS1_SFF_71_Q_reg ( .D(
        Inst_forkAE_CipherInst_RF_RS1_SFF_71_N3), .SI(1'b0), .SE(1'b0), .CK(
        clk), .SN(1'b1), .Q(Inst_forkAE_CipherInst_RF_S_MID_D1[71]) );
  SDFFSQX2 Inst_forkAE_ControlInst_fsm_state_reg_1_ ( .D(
        Inst_forkAE_ControlInst_n32), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_ControlInst_fsm_state_1_) );
  AND2X2 U1 ( .A(Inst_forkAE_ControlInst_fsm_state_1_), .B(n2244), .Y(n1) );
  AND2X2 U2 ( .A(a_data), .B(n145), .Y(n5) );
  AND2X2 U3 ( .A(n1989), .B(n145), .Y(n7) );
  NAND2X2 U4 ( .A(n2244), .B(Inst_forkAE_CipherInst_CL_n34), .Y(n2005) );
  NAND2X2 U5 ( .A(dec), .B(n245), .Y(n2244) );
  INVX2 U6 ( .A(n2244), .Y(n1989) );
  INVX2 U7 ( .A(n2255), .Y(n2312) );
  INVX2 U8 ( .A(n2722), .Y(n2258) );
  NAND2X1 U9 ( .A(n2293), .B(n310), .Y(n2722) );
  INVX2 U10 ( .A(n2274), .Y(n2293) );
  NOR2X4 U11 ( .A(n145), .B(n2244), .Y(n5443) );
  CLKNAND2X4 U12 ( .A(n1989), .B(n2267), .Y(n2274) );
  NAND2X3 U13 ( .A(Inst_forkAE_CipherInst_LAST), .B(n1989), .Y(n2267) );
  NAND2X4 U14 ( .A(Inst_forkAE_CipherInst_LAST), .B(n2244), .Y(n2273) );
  NAND2X4 U15 ( .A(Block_Size[0]), .B(n3977), .Y(n2288) );
  NAND3X2 U16 ( .A(n255), .B(n159), .C(n2000), .Y(n2302) );
  BUFX2 U17 ( .A(n380), .Y(n371) );
  BUFX2 U18 ( .A(n378), .Y(n376) );
  BUFX2 U19 ( .A(n378), .Y(n375) );
  BUFX2 U20 ( .A(n379), .Y(n374) );
  BUFX2 U21 ( .A(n379), .Y(n373) );
  BUFX2 U22 ( .A(n379), .Y(n372) );
  BUFX2 U23 ( .A(n380), .Y(n370) );
  BUFX2 U24 ( .A(n385), .Y(n355) );
  BUFX2 U25 ( .A(n385), .Y(n356) );
  BUFX2 U26 ( .A(n382), .Y(n363) );
  BUFX2 U27 ( .A(n384), .Y(n357) );
  BUFX2 U28 ( .A(n384), .Y(n358) );
  BUFX2 U29 ( .A(n384), .Y(n359) );
  BUFX2 U30 ( .A(n383), .Y(n360) );
  BUFX2 U31 ( .A(n383), .Y(n361) );
  BUFX2 U32 ( .A(n383), .Y(n362) );
  BUFX2 U33 ( .A(n382), .Y(n364) );
  BUFX2 U34 ( .A(n382), .Y(n365) );
  BUFX2 U35 ( .A(n381), .Y(n366) );
  BUFX2 U36 ( .A(n381), .Y(n367) );
  BUFX2 U37 ( .A(n381), .Y(n368) );
  BUFX2 U38 ( .A(n380), .Y(n369) );
  BUFX2 U39 ( .A(n378), .Y(n377) );
  INVX2 U40 ( .A(n412), .Y(n409) );
  BUFX2 U41 ( .A(n241), .Y(n222) );
  BUFX2 U42 ( .A(n241), .Y(n223) );
  BUFX2 U43 ( .A(n241), .Y(n224) );
  BUFX2 U44 ( .A(n240), .Y(n225) );
  BUFX2 U45 ( .A(n240), .Y(n226) );
  BUFX2 U46 ( .A(n242), .Y(n220) );
  BUFX2 U47 ( .A(n242), .Y(n221) );
  BUFX2 U48 ( .A(n239), .Y(n230) );
  BUFX2 U49 ( .A(n238), .Y(n231) );
  BUFX2 U50 ( .A(n238), .Y(n232) );
  BUFX2 U51 ( .A(n238), .Y(n233) );
  BUFX2 U52 ( .A(n237), .Y(n234) );
  BUFX2 U53 ( .A(n237), .Y(n235) );
  BUFX2 U54 ( .A(n240), .Y(n227) );
  BUFX2 U55 ( .A(n239), .Y(n228) );
  BUFX2 U56 ( .A(n239), .Y(n229) );
  BUFX2 U57 ( .A(n242), .Y(n219) );
  INVX2 U58 ( .A(n412), .Y(n410) );
  INVX2 U59 ( .A(n413), .Y(n408) );
  BUFX2 U60 ( .A(n214), .Y(n193) );
  BUFX2 U61 ( .A(n213), .Y(n194) );
  BUFX2 U62 ( .A(n213), .Y(n195) );
  BUFX2 U63 ( .A(n213), .Y(n196) );
  BUFX2 U64 ( .A(n212), .Y(n197) );
  BUFX2 U65 ( .A(n212), .Y(n198) );
  BUFX2 U66 ( .A(n214), .Y(n191) );
  BUFX2 U67 ( .A(n214), .Y(n192) );
  BUFX2 U68 ( .A(n211), .Y(n202) );
  BUFX2 U69 ( .A(n210), .Y(n203) );
  BUFX2 U70 ( .A(n210), .Y(n204) );
  BUFX2 U71 ( .A(n210), .Y(n205) );
  BUFX2 U72 ( .A(n212), .Y(n199) );
  BUFX2 U73 ( .A(n211), .Y(n200) );
  BUFX2 U74 ( .A(n211), .Y(n201) );
  BUFX2 U75 ( .A(n237), .Y(n236) );
  BUFX2 U76 ( .A(n415), .Y(n412) );
  BUFX2 U77 ( .A(n415), .Y(n413) );
  BUFX2 U78 ( .A(n415), .Y(n414) );
  BUFX2 U79 ( .A(n387), .Y(n381) );
  BUFX2 U80 ( .A(n387), .Y(n380) );
  BUFX2 U81 ( .A(n387), .Y(n382) );
  BUFX2 U82 ( .A(n386), .Y(n384) );
  BUFX2 U83 ( .A(n386), .Y(n383) );
  BUFX2 U84 ( .A(n388), .Y(n378) );
  BUFX2 U85 ( .A(n388), .Y(n379) );
  BUFX2 U86 ( .A(n216), .Y(n213) );
  BUFX2 U87 ( .A(n216), .Y(n214) );
  BUFX2 U88 ( .A(n217), .Y(n210) );
  BUFX2 U89 ( .A(n217), .Y(n212) );
  BUFX2 U90 ( .A(n217), .Y(n211) );
  BUFX2 U91 ( .A(n243), .Y(n241) );
  BUFX2 U92 ( .A(n244), .Y(n238) );
  BUFX2 U93 ( .A(n244), .Y(n237) );
  BUFX2 U94 ( .A(n243), .Y(n240) );
  BUFX2 U95 ( .A(n244), .Y(n239) );
  BUFX2 U96 ( .A(n243), .Y(n242) );
  BUFX2 U97 ( .A(n142), .Y(n123) );
  BUFX2 U98 ( .A(n140), .Y(n130) );
  BUFX2 U99 ( .A(n139), .Y(n132) );
  BUFX2 U100 ( .A(n139), .Y(n133) );
  BUFX2 U101 ( .A(n139), .Y(n134) );
  BUFX2 U102 ( .A(n138), .Y(n135) );
  BUFX2 U103 ( .A(n138), .Y(n136) );
  BUFX2 U104 ( .A(n138), .Y(n137) );
  BUFX2 U105 ( .A(n140), .Y(n131) );
  BUFX2 U106 ( .A(n142), .Y(n124) );
  BUFX2 U107 ( .A(n142), .Y(n125) );
  BUFX2 U108 ( .A(n141), .Y(n128) );
  BUFX2 U109 ( .A(n141), .Y(n127) );
  BUFX2 U110 ( .A(n141), .Y(n126) );
  BUFX2 U111 ( .A(n140), .Y(n129) );
  BUFX2 U112 ( .A(n386), .Y(n385) );
  BUFX2 U113 ( .A(n404), .Y(n398) );
  BUFX2 U114 ( .A(n404), .Y(n397) );
  BUFX2 U115 ( .A(n403), .Y(n400) );
  BUFX2 U116 ( .A(n403), .Y(n401) );
  BUFX2 U117 ( .A(n305), .Y(n296) );
  BUFX2 U118 ( .A(n304), .Y(n297) );
  BUFX2 U119 ( .A(n304), .Y(n299) );
  BUFX2 U120 ( .A(n405), .Y(n395) );
  BUFX2 U121 ( .A(n404), .Y(n399) );
  BUFX2 U122 ( .A(n405), .Y(n396) );
  BUFX2 U123 ( .A(n406), .Y(n393) );
  BUFX2 U124 ( .A(n406), .Y(n392) );
  BUFX2 U125 ( .A(n406), .Y(n391) );
  BUFX2 U126 ( .A(n405), .Y(n394) );
  BUFX2 U127 ( .A(n407), .Y(n390) );
  BUFX2 U128 ( .A(n407), .Y(n389) );
  BUFX2 U129 ( .A(n304), .Y(n298) );
  BUFX2 U130 ( .A(n305), .Y(n295) );
  BUFX2 U131 ( .A(n303), .Y(n301) );
  BUFX2 U132 ( .A(n303), .Y(n300) );
  BUFX2 U133 ( .A(n305), .Y(n294) );
  BUFX2 U134 ( .A(n271), .Y(n266) );
  BUFX2 U135 ( .A(n271), .Y(n265) );
  BUFX2 U136 ( .A(n270), .Y(n267) );
  BUFX2 U137 ( .A(n272), .Y(n261) );
  BUFX2 U138 ( .A(n270), .Y(n268) );
  BUFX2 U139 ( .A(n272), .Y(n263) );
  BUFX2 U140 ( .A(n272), .Y(n262) );
  BUFX2 U141 ( .A(n403), .Y(n402) );
  BUFX2 U142 ( .A(n271), .Y(n264) );
  BUFX2 U143 ( .A(n215), .Y(n190) );
  BUFX2 U144 ( .A(n216), .Y(n215) );
  BUFX2 U145 ( .A(n209), .Y(n206) );
  BUFX2 U146 ( .A(n209), .Y(n207) );
  INVX2 U147 ( .A(n289), .Y(n276) );
  INVX2 U148 ( .A(n289), .Y(n277) );
  INVX2 U149 ( .A(n288), .Y(n278) );
  INVX2 U150 ( .A(n288), .Y(n279) );
  INVX2 U151 ( .A(n288), .Y(n280) );
  INVX2 U152 ( .A(n287), .Y(n281) );
  INVX2 U153 ( .A(n287), .Y(n282) );
  INVX2 U154 ( .A(n287), .Y(n283) );
  INVX2 U155 ( .A(n290), .Y(n275) );
  INVX2 U156 ( .A(n291), .Y(n274) );
  BUFX2 U157 ( .A(n209), .Y(n208) );
  BUFX2 U158 ( .A(n270), .Y(n269) );
  BUFX2 U159 ( .A(n303), .Y(n302) );
  BUFX2 U160 ( .A(n293), .Y(n287) );
  BUFX2 U161 ( .A(n293), .Y(n290) );
  BUFX2 U162 ( .A(n293), .Y(n288) );
  BUFX2 U163 ( .A(n286), .Y(n289) );
  BUFX2 U164 ( .A(n293), .Y(n291) );
  BUFX2 U165 ( .A(n2260), .Y(n272) );
  BUFX2 U166 ( .A(n2260), .Y(n270) );
  BUFX2 U167 ( .A(n2260), .Y(n271) );
  BUFX2 U168 ( .A(n4963), .Y(n387) );
  BUFX2 U169 ( .A(n4963), .Y(n386) );
  BUFX2 U170 ( .A(n416), .Y(n411) );
  BUFX2 U171 ( .A(n7), .Y(n416) );
  BUFX2 U172 ( .A(n5192), .Y(n403) );
  BUFX2 U173 ( .A(n5192), .Y(n406) );
  BUFX2 U174 ( .A(n5192), .Y(n404) );
  BUFX2 U175 ( .A(n5192), .Y(n405) );
  BUFX2 U176 ( .A(n4963), .Y(n388) );
  BUFX2 U177 ( .A(n2286), .Y(n304) );
  BUFX2 U178 ( .A(n2286), .Y(n305) );
  BUFX2 U179 ( .A(n2286), .Y(n303) );
  BUFX2 U180 ( .A(n5192), .Y(n407) );
  BUFX2 U181 ( .A(n2249), .Y(n244) );
  BUFX2 U182 ( .A(n2249), .Y(n243) );
  BUFX2 U183 ( .A(n2248), .Y(n217) );
  BUFX2 U184 ( .A(n2248), .Y(n216) );
  BUFX2 U185 ( .A(n293), .Y(n292) );
  BUFX2 U186 ( .A(n456), .Y(n417) );
  BUFX2 U187 ( .A(n454), .Y(n424) );
  BUFX2 U188 ( .A(n455), .Y(n421) );
  BUFX2 U189 ( .A(n455), .Y(n422) );
  BUFX2 U190 ( .A(n454), .Y(n423) );
  BUFX2 U191 ( .A(n454), .Y(n425) );
  BUFX2 U192 ( .A(n456), .Y(n418) );
  BUFX2 U193 ( .A(n456), .Y(n419) );
  BUFX2 U194 ( .A(n455), .Y(n420) );
  BUFX2 U195 ( .A(n453), .Y(n426) );
  BUFX2 U196 ( .A(n451), .Y(n434) );
  BUFX2 U197 ( .A(n453), .Y(n427) );
  BUFX2 U198 ( .A(n453), .Y(n428) );
  BUFX2 U199 ( .A(n451), .Y(n433) );
  BUFX2 U200 ( .A(n452), .Y(n430) );
  BUFX2 U201 ( .A(n452), .Y(n431) );
  BUFX2 U202 ( .A(n450), .Y(n435) );
  BUFX2 U203 ( .A(n452), .Y(n429) );
  BUFX2 U204 ( .A(n451), .Y(n432) );
  BUFX2 U205 ( .A(n450), .Y(n436) );
  BUFX2 U206 ( .A(n450), .Y(n437) );
  BUFX2 U207 ( .A(n448), .Y(n443) );
  BUFX2 U208 ( .A(n449), .Y(n440) );
  BUFX2 U209 ( .A(n448), .Y(n441) );
  BUFX2 U210 ( .A(n449), .Y(n439) );
  BUFX2 U211 ( .A(n449), .Y(n438) );
  BUFX2 U212 ( .A(n448), .Y(n442) );
  BUFX2 U213 ( .A(n7), .Y(n415) );
  BUFX2 U214 ( .A(n143), .Y(n142) );
  BUFX2 U215 ( .A(n143), .Y(n141) );
  BUFX2 U216 ( .A(n143), .Y(n140) );
  BUFX2 U217 ( .A(n218), .Y(n209) );
  BUFX2 U218 ( .A(n2248), .Y(n218) );
  BUFX2 U219 ( .A(n144), .Y(n139) );
  BUFX2 U220 ( .A(n144), .Y(n138) );
  BUFX2 U221 ( .A(n60), .Y(n14) );
  BUFX2 U222 ( .A(n60), .Y(n15) );
  BUFX2 U223 ( .A(n57), .Y(n23) );
  BUFX2 U224 ( .A(n57), .Y(n24) );
  BUFX2 U225 ( .A(n56), .Y(n25) );
  BUFX2 U226 ( .A(n56), .Y(n26) );
  BUFX2 U227 ( .A(n56), .Y(n27) );
  BUFX2 U228 ( .A(n55), .Y(n28) );
  BUFX2 U229 ( .A(n55), .Y(n30) );
  BUFX2 U230 ( .A(n55), .Y(n29) );
  BUFX2 U231 ( .A(n59), .Y(n16) );
  BUFX2 U232 ( .A(n59), .Y(n17) );
  BUFX2 U233 ( .A(n59), .Y(n18) );
  BUFX2 U234 ( .A(n58), .Y(n19) );
  BUFX2 U235 ( .A(n58), .Y(n20) );
  BUFX2 U236 ( .A(n58), .Y(n21) );
  BUFX2 U237 ( .A(n57), .Y(n22) );
  BUFX2 U238 ( .A(n53), .Y(n34) );
  INVX2 U239 ( .A(n321), .Y(n316) );
  INVX2 U240 ( .A(n321), .Y(n315) );
  INVX2 U241 ( .A(n317), .Y(n308) );
  INVX2 U242 ( .A(n318), .Y(n310) );
  INVX2 U243 ( .A(n318), .Y(n309) );
  INVX2 U244 ( .A(n320), .Y(n312) );
  INVX2 U245 ( .A(n321), .Y(n314) );
  INVX2 U246 ( .A(n320), .Y(n313) );
  INVX2 U247 ( .A(n317), .Y(n307) );
  INVX2 U248 ( .A(n317), .Y(n306) );
  INVX2 U249 ( .A(n318), .Y(n311) );
  BUFX2 U250 ( .A(n54), .Y(n31) );
  BUFX2 U251 ( .A(n53), .Y(n35) );
  BUFX2 U252 ( .A(n54), .Y(n32) );
  BUFX2 U253 ( .A(n51), .Y(n40) );
  BUFX2 U254 ( .A(n52), .Y(n39) );
  BUFX2 U255 ( .A(n52), .Y(n38) );
  BUFX2 U256 ( .A(n52), .Y(n37) );
  BUFX2 U257 ( .A(n53), .Y(n36) );
  BUFX2 U258 ( .A(n49), .Y(n47) );
  BUFX2 U259 ( .A(n49), .Y(n46) );
  BUFX2 U260 ( .A(n50), .Y(n45) );
  BUFX2 U261 ( .A(n50), .Y(n44) );
  BUFX2 U262 ( .A(n50), .Y(n43) );
  BUFX2 U263 ( .A(n51), .Y(n42) );
  BUFX2 U264 ( .A(n51), .Y(n41) );
  BUFX2 U265 ( .A(n54), .Y(n33) );
  BUFX2 U266 ( .A(n259), .Y(n245) );
  BUFX2 U267 ( .A(n258), .Y(n247) );
  BUFX2 U268 ( .A(n258), .Y(n248) );
  BUFX2 U269 ( .A(n257), .Y(n252) );
  BUFX2 U270 ( .A(n257), .Y(n251) );
  BUFX2 U271 ( .A(n257), .Y(n250) );
  BUFX2 U272 ( .A(n258), .Y(n249) );
  BUFX2 U273 ( .A(n256), .Y(n253) );
  BUFX2 U274 ( .A(n259), .Y(n246) );
  BUFX2 U275 ( .A(n256), .Y(n254) );
  BUFX2 U276 ( .A(n91), .Y(n65) );
  BUFX2 U277 ( .A(n91), .Y(n66) );
  BUFX2 U278 ( .A(n88), .Y(n74) );
  BUFX2 U279 ( .A(n88), .Y(n75) );
  BUFX2 U280 ( .A(n87), .Y(n76) );
  BUFX2 U281 ( .A(n87), .Y(n77) );
  BUFX2 U282 ( .A(n87), .Y(n78) );
  BUFX2 U283 ( .A(n86), .Y(n79) );
  BUFX2 U284 ( .A(n86), .Y(n80) );
  BUFX2 U285 ( .A(n86), .Y(n81) );
  BUFX2 U286 ( .A(n88), .Y(n73) );
  BUFX2 U287 ( .A(n89), .Y(n72) );
  BUFX2 U288 ( .A(n89), .Y(n71) );
  BUFX2 U289 ( .A(n89), .Y(n70) );
  BUFX2 U290 ( .A(n90), .Y(n69) );
  BUFX2 U291 ( .A(n90), .Y(n68) );
  BUFX2 U292 ( .A(n90), .Y(n67) );
  BUFX2 U293 ( .A(n121), .Y(n98) );
  BUFX2 U294 ( .A(n121), .Y(n99) );
  BUFX2 U295 ( .A(n121), .Y(n100) );
  BUFX2 U296 ( .A(n120), .Y(n101) );
  BUFX2 U297 ( .A(n120), .Y(n102) );
  BUFX2 U298 ( .A(n118), .Y(n107) );
  BUFX2 U299 ( .A(n119), .Y(n105) );
  BUFX2 U300 ( .A(n119), .Y(n106) );
  BUFX2 U301 ( .A(n119), .Y(n104) );
  BUFX2 U302 ( .A(n120), .Y(n103) );
  BUFX2 U303 ( .A(n122), .Y(n97) );
  BUFX2 U304 ( .A(n122), .Y(n96) );
  BUFX2 U305 ( .A(n118), .Y(n108) );
  BUFX2 U306 ( .A(n116), .Y(n114) );
  BUFX2 U307 ( .A(n116), .Y(n113) );
  BUFX2 U308 ( .A(n117), .Y(n112) );
  BUFX2 U309 ( .A(n117), .Y(n111) );
  BUFX2 U310 ( .A(n118), .Y(n109) );
  BUFX2 U311 ( .A(n117), .Y(n110) );
  BUFX2 U312 ( .A(n273), .Y(n260) );
  BUFX2 U313 ( .A(n2260), .Y(n273) );
  INVX2 U314 ( .A(n353), .Y(n325) );
  INVX2 U315 ( .A(n353), .Y(n326) );
  INVX2 U316 ( .A(n352), .Y(n327) );
  INVX2 U317 ( .A(n351), .Y(n330) );
  INVX2 U318 ( .A(n351), .Y(n331) );
  INVX2 U319 ( .A(n350), .Y(n334) );
  INVX2 U320 ( .A(n350), .Y(n333) );
  INVX2 U321 ( .A(n351), .Y(n332) );
  INVX2 U322 ( .A(n350), .Y(n335) );
  INVX2 U323 ( .A(n352), .Y(n329) );
  INVX2 U324 ( .A(n352), .Y(n328) );
  INVX2 U325 ( .A(n349), .Y(n336) );
  INVX2 U326 ( .A(n347), .Y(n344) );
  INVX2 U327 ( .A(n347), .Y(n343) );
  INVX2 U328 ( .A(n347), .Y(n342) );
  INVX2 U329 ( .A(n348), .Y(n341) );
  INVX2 U330 ( .A(n349), .Y(n338) );
  INVX2 U331 ( .A(n348), .Y(n339) );
  INVX2 U332 ( .A(n349), .Y(n337) );
  INVX2 U333 ( .A(n348), .Y(n340) );
  INVX2 U334 ( .A(n286), .Y(n285) );
  INVX2 U335 ( .A(n346), .Y(n345) );
  INVX2 U336 ( .A(n286), .Y(n284) );
  INVX2 U337 ( .A(n183), .Y(n171) );
  INVX2 U338 ( .A(n183), .Y(n172) );
  INVX2 U339 ( .A(n182), .Y(n176) );
  INVX2 U340 ( .A(n181), .Y(n177) );
  INVX2 U341 ( .A(n181), .Y(n178) );
  INVX2 U342 ( .A(n181), .Y(n179) );
  INVX2 U343 ( .A(n183), .Y(n173) );
  INVX2 U344 ( .A(n182), .Y(n174) );
  INVX2 U345 ( .A(n182), .Y(n175) );
  INVX2 U346 ( .A(n185), .Y(n167) );
  INVX2 U347 ( .A(n184), .Y(n168) );
  INVX2 U348 ( .A(n184), .Y(n169) );
  INVX2 U349 ( .A(n184), .Y(n170) );
  INVX2 U350 ( .A(n185), .Y(n166) );
  BUFX2 U351 ( .A(n49), .Y(n48) );
  BUFX2 U352 ( .A(n256), .Y(n255) );
  INVX2 U353 ( .A(n186), .Y(n165) );
  BUFX2 U354 ( .A(n116), .Y(n115) );
  BUFX2 U355 ( .A(n2254), .Y(n257) );
  BUFX2 U356 ( .A(n2254), .Y(n258) );
  BUFX2 U357 ( .A(n2254), .Y(n256) );
  BUFX2 U358 ( .A(n1), .Y(n347) );
  BUFX2 U359 ( .A(n1), .Y(n346) );
  BUFX2 U360 ( .A(n1), .Y(n349) );
  BUFX2 U361 ( .A(n1), .Y(n348) );
  BUFX2 U362 ( .A(n1), .Y(n351) );
  BUFX2 U363 ( .A(n1), .Y(n350) );
  BUFX2 U364 ( .A(n1), .Y(n352) );
  BUFX2 U365 ( .A(n293), .Y(n286) );
  INVX2 U366 ( .A(n2266), .Y(n293) );
  BUFX2 U367 ( .A(n350), .Y(n353) );
  BUFX2 U368 ( .A(n324), .Y(n318) );
  BUFX2 U369 ( .A(n324), .Y(n317) );
  BUFX2 U370 ( .A(n323), .Y(n320) );
  BUFX2 U371 ( .A(n324), .Y(n319) );
  BUFX2 U372 ( .A(n323), .Y(n321) );
  BUFX2 U373 ( .A(n188), .Y(n181) );
  BUFX2 U374 ( .A(n188), .Y(n183) );
  BUFX2 U375 ( .A(n188), .Y(n182) );
  BUFX2 U376 ( .A(n187), .Y(n184) );
  BUFX2 U377 ( .A(n187), .Y(n185) );
  BUFX2 U378 ( .A(n1069), .Y(n121) );
  BUFX2 U379 ( .A(n1069), .Y(n116) );
  BUFX2 U380 ( .A(n1069), .Y(n119) );
  BUFX2 U381 ( .A(n1069), .Y(n118) );
  BUFX2 U382 ( .A(n1069), .Y(n120) );
  BUFX2 U383 ( .A(n1069), .Y(n117) );
  BUFX2 U384 ( .A(n2254), .Y(n259) );
  BUFX2 U385 ( .A(n1069), .Y(n122) );
  BUFX2 U386 ( .A(n1071), .Y(n143) );
  BUFX2 U387 ( .A(n1071), .Y(n144) );
  BUFX2 U388 ( .A(n349), .Y(n354) );
  BUFX2 U389 ( .A(n187), .Y(n186) );
  BUFX2 U390 ( .A(n447), .Y(n444) );
  BUFX2 U391 ( .A(n447), .Y(n445) );
  BUFX2 U392 ( .A(n62), .Y(n56) );
  BUFX2 U393 ( .A(n63), .Y(n52) );
  BUFX2 U394 ( .A(n62), .Y(n55) );
  BUFX2 U395 ( .A(n64), .Y(n49) );
  BUFX2 U396 ( .A(n61), .Y(n59) );
  BUFX2 U397 ( .A(n64), .Y(n50) );
  BUFX2 U398 ( .A(n61), .Y(n58) );
  BUFX2 U399 ( .A(n62), .Y(n57) );
  BUFX2 U400 ( .A(n63), .Y(n53) );
  BUFX2 U401 ( .A(n64), .Y(n51) );
  BUFX2 U402 ( .A(n63), .Y(n54) );
  BUFX2 U403 ( .A(n457), .Y(n454) );
  BUFX2 U404 ( .A(n457), .Y(n456) );
  BUFX2 U405 ( .A(n457), .Y(n455) );
  BUFX2 U406 ( .A(n458), .Y(n453) );
  BUFX2 U407 ( .A(n458), .Y(n452) );
  BUFX2 U408 ( .A(n458), .Y(n451) );
  BUFX2 U409 ( .A(n459), .Y(n450) );
  BUFX2 U410 ( .A(n459), .Y(n449) );
  BUFX2 U411 ( .A(n459), .Y(n448) );
  BUFX2 U412 ( .A(n93), .Y(n87) );
  BUFX2 U413 ( .A(n93), .Y(n86) );
  BUFX2 U414 ( .A(n93), .Y(n88) );
  BUFX2 U415 ( .A(n92), .Y(n89) );
  BUFX2 U416 ( .A(n92), .Y(n90) );
  BUFX2 U417 ( .A(n164), .Y(n145) );
  BUFX2 U418 ( .A(n160), .Y(n159) );
  BUFX2 U419 ( .A(n161), .Y(n155) );
  BUFX2 U420 ( .A(n160), .Y(n157) );
  BUFX2 U421 ( .A(n160), .Y(n158) );
  BUFX2 U422 ( .A(n162), .Y(n153) );
  BUFX2 U423 ( .A(n161), .Y(n156) );
  BUFX2 U424 ( .A(n161), .Y(n154) );
  BUFX2 U425 ( .A(n163), .Y(n148) );
  BUFX2 U426 ( .A(n163), .Y(n149) );
  BUFX2 U427 ( .A(n163), .Y(n150) );
  BUFX2 U428 ( .A(n162), .Y(n151) );
  BUFX2 U429 ( .A(n164), .Y(n146) );
  BUFX2 U430 ( .A(n164), .Y(n147) );
  BUFX2 U431 ( .A(n162), .Y(n152) );
  BUFX2 U432 ( .A(n85), .Y(n82) );
  BUFX2 U433 ( .A(n85), .Y(n83) );
  BUFX2 U434 ( .A(n92), .Y(n91) );
  BUFX2 U435 ( .A(n61), .Y(n60) );
  BUFX2 U436 ( .A(n447), .Y(n446) );
  BUFX2 U437 ( .A(n85), .Y(n84) );
  BUFX2 U438 ( .A(n323), .Y(n322) );
  OAI2B11X2 U439 ( .A1N(n286), .A0(n3732), .B0(n4165), .C0(n4166), .Y(n4164)
         );
  BUFX2 U440 ( .A(Inst_forkAE_CipherInst_KE_CLK_K), .Y(n457) );
  BUFX2 U441 ( .A(Inst_forkAE_CipherInst_KE_CLK_K), .Y(n458) );
  BUFX2 U442 ( .A(Inst_forkAE_CipherInst_KE_CLK_K), .Y(n459) );
  BUFX2 U443 ( .A(n587), .Y(n61) );
  BUFX2 U444 ( .A(n587), .Y(n62) );
  BUFX2 U445 ( .A(n587), .Y(n64) );
  BUFX2 U446 ( .A(n587), .Y(n63) );
  BUFX2 U447 ( .A(n189), .Y(n180) );
  BUFX2 U448 ( .A(n5), .Y(n189) );
  BUFX2 U449 ( .A(n1985), .Y(n160) );
  BUFX2 U450 ( .A(n1985), .Y(n161) );
  BUFX2 U451 ( .A(n1985), .Y(n163) );
  BUFX2 U452 ( .A(n1985), .Y(n164) );
  BUFX2 U453 ( .A(n1985), .Y(n162) );
  BUFX2 U454 ( .A(n8), .Y(n324) );
  BUFX2 U455 ( .A(n8), .Y(n323) );
  BUFX2 U456 ( .A(n94), .Y(n85) );
  BUFX2 U457 ( .A(n95), .Y(n94) );
  BUFX2 U458 ( .A(n5), .Y(n188) );
  BUFX2 U459 ( .A(n5), .Y(n187) );
  BUFX2 U460 ( .A(n95), .Y(n93) );
  BUFX2 U461 ( .A(n95), .Y(n92) );
  BUFX2 U462 ( .A(n460), .Y(n447) );
  BUFX2 U463 ( .A(Inst_forkAE_CipherInst_KE_CLK_K), .Y(n460) );
  OR3X2 U464 ( .A(Inst_forkAE_CipherInst_CL_COUNTER_0_), .B(
        Inst_forkAE_CipherInst_CL_COUNTER_2_), .C(n2), .Y(n8) );
  BUFX2 U465 ( .A(n588), .Y(n95) );
  CLKNAND2X2 U466 ( .A(n485), .B(n5715), .Y(n5716) );
  MXI2X1 U467 ( .A(Inst_forkAE_CipherInst_TK1_DEC_48_), .B(n3), .S0(done), .Y(
        n485) );
  XOR2X1 U468 ( .A(Inst_forkAE_CipherInst_CL_COUNTER_0_), .B(n2), .Y(n5719) );
  CLKINVX1 U469 ( .A(n486), .Y(Tag2[9]) );
  CLKINVX1 U470 ( .A(n487), .Y(Tag2[97]) );
  CLKINVX1 U471 ( .A(n488), .Y(Tag2[96]) );
  CLKINVX1 U472 ( .A(n489), .Y(Tag2[95]) );
  CLKINVX1 U473 ( .A(n490), .Y(Tag2[93]) );
  CLKINVX1 U474 ( .A(n491), .Y(Tag2[90]) );
  CLKINVX1 U475 ( .A(n492), .Y(Tag2[87]) );
  CLKINVX1 U476 ( .A(n493), .Y(Tag2[85]) );
  CLKINVX1 U477 ( .A(n494), .Y(Tag2[82]) );
  CLKINVX1 U478 ( .A(n495), .Y(Tag2[77]) );
  CLKINVX1 U479 ( .A(n496), .Y(Tag2[74]) );
  CLKINVX1 U480 ( .A(n497), .Y(Tag2[6]) );
  CLKINVX1 U481 ( .A(n498), .Y(Tag2[69]) );
  CLKINVX1 U482 ( .A(n499), .Y(Tag2[66]) );
  CLKINVX1 U483 ( .A(n500), .Y(Tag2[62]) );
  CLKINVX1 U484 ( .A(n501), .Y(Tag2[61]) );
  CLKINVX1 U485 ( .A(n502), .Y(Tag2[57]) );
  CLKINVX1 U486 ( .A(n503), .Y(Tag2[54]) );
  CLKINVX1 U487 ( .A(n504), .Y(Tag2[53]) );
  CLKINVX1 U488 ( .A(n505), .Y(Tag2[49]) );
  CLKINVX1 U489 ( .A(n506), .Y(Tag2[46]) );
  CLKINVX1 U490 ( .A(n507), .Y(Tag2[45]) );
  CLKINVX1 U491 ( .A(n508), .Y(Tag2[41]) );
  CLKINVX1 U492 ( .A(n509), .Y(Tag2[38]) );
  CLKINVX1 U493 ( .A(n510), .Y(Tag2[37]) );
  CLKINVX1 U494 ( .A(n511), .Y(Tag2[33]) );
  CLKINVX1 U495 ( .A(n512), .Y(Tag2[30]) );
  CLKINVX1 U496 ( .A(n513), .Y(Tag2[25]) );
  CLKINVX1 U497 ( .A(n514), .Y(Tag2[22]) );
  CLKINVX1 U498 ( .A(n515), .Y(Tag2[1]) );
  CLKINVX1 U499 ( .A(n516), .Y(Tag2[14]) );
  CLKINVX1 U500 ( .A(n517), .Y(Tag2[126]) );
  CLKINVX1 U501 ( .A(n518), .Y(Tag2[125]) );
  CLKINVX1 U502 ( .A(n519), .Y(Tag2[121]) );
  CLKINVX1 U503 ( .A(n520), .Y(Tag2[118]) );
  CLKINVX1 U504 ( .A(n521), .Y(Tag2[117]) );
  CLKINVX1 U505 ( .A(n522), .Y(Tag2[113]) );
  CLKINVX1 U506 ( .A(n523), .Y(Tag2[110]) );
  CLKINVX1 U507 ( .A(n524), .Y(Tag2[109]) );
  CLKINVX1 U508 ( .A(n525), .Y(Tag2[105]) );
  CLKINVX1 U509 ( .A(n526), .Y(Tag2[102]) );
  CLKINVX1 U510 ( .A(n527), .Y(Tag2[101]) );
  CLKINVX1 U511 ( .A(n528), .Y(Tag1[97]) );
  CLKINVX1 U512 ( .A(n529), .Y(Tag1[96]) );
  CLKINVX1 U513 ( .A(n530), .Y(Tag1[94]) );
  CLKINVX1 U514 ( .A(n531), .Y(Tag1[89]) );
  CLKINVX1 U515 ( .A(n532), .Y(Tag1[86]) );
  CLKINVX1 U516 ( .A(n533), .Y(Tag1[81]) );
  CLKINVX1 U517 ( .A(n534), .Y(Tag1[78]) );
  CLKINVX1 U518 ( .A(n535), .Y(Tag1[73]) );
  CLKINVX1 U519 ( .A(n536), .Y(Tag1[70]) );
  CLKINVX1 U520 ( .A(n537), .Y(Tag1[6]) );
  CLKINVX1 U521 ( .A(n538), .Y(Tag1[65]) );
  CLKINVX1 U522 ( .A(n539), .Y(Tag1[62]) );
  CLKINVX1 U523 ( .A(n540), .Y(Tag1[61]) );
  CLKINVX1 U524 ( .A(n541), .Y(Tag1[60]) );
  CLKINVX1 U525 ( .A(n542), .Y(Tag1[57]) );
  CLKINVX1 U526 ( .A(n543), .Y(Tag1[56]) );
  CLKINVX1 U527 ( .A(n544), .Y(Tag1[54]) );
  CLKINVX1 U528 ( .A(n545), .Y(Tag1[53]) );
  CLKINVX1 U529 ( .A(n546), .Y(Tag1[52]) );
  CLKINVX1 U530 ( .A(n547), .Y(Tag1[49]) );
  CLKINVX1 U531 ( .A(n548), .Y(Tag1[48]) );
  CLKINVX1 U532 ( .A(n549), .Y(Tag1[46]) );
  CLKINVX1 U533 ( .A(n550), .Y(Tag1[45]) );
  CLKINVX1 U534 ( .A(n551), .Y(Tag1[44]) );
  CLKINVX1 U535 ( .A(n552), .Y(Tag1[41]) );
  CLKINVX1 U536 ( .A(n553), .Y(Tag1[40]) );
  CLKINVX1 U537 ( .A(n554), .Y(Tag1[38]) );
  CLKINVX1 U538 ( .A(n555), .Y(Tag1[37]) );
  CLKINVX1 U539 ( .A(n556), .Y(Tag1[36]) );
  CLKINVX1 U540 ( .A(n557), .Y(Tag1[33]) );
  CLKINVX1 U541 ( .A(n558), .Y(Tag1[32]) );
  CLKINVX1 U542 ( .A(n559), .Y(Tag1[30]) );
  CLKINVX1 U543 ( .A(n560), .Y(Tag1[22]) );
  CLKINVX1 U544 ( .A(n561), .Y(Tag1[21]) );
  CLKINVX1 U545 ( .A(n562), .Y(Tag1[1]) );
  CLKINVX1 U546 ( .A(n563), .Y(Tag1[17]) );
  CLKINVX1 U547 ( .A(n564), .Y(Tag1[14]) );
  CLKINVX1 U548 ( .A(n565), .Y(Tag1[13]) );
  CLKINVX1 U549 ( .A(n566), .Y(Tag1[126]) );
  CLKINVX1 U550 ( .A(n567), .Y(Tag1[125]) );
  CLKINVX1 U551 ( .A(n568), .Y(Tag1[124]) );
  CLKINVX1 U552 ( .A(n569), .Y(Tag1[121]) );
  CLKINVX1 U553 ( .A(n570), .Y(Tag1[120]) );
  CLKINVX1 U554 ( .A(n571), .Y(Tag1[118]) );
  CLKINVX1 U555 ( .A(n572), .Y(Tag1[117]) );
  CLKINVX1 U556 ( .A(n573), .Y(Tag1[116]) );
  CLKINVX1 U557 ( .A(n574), .Y(Tag1[113]) );
  CLKINVX1 U558 ( .A(n575), .Y(Tag1[112]) );
  CLKINVX1 U559 ( .A(n576), .Y(Tag1[110]) );
  CLKINVX1 U560 ( .A(n577), .Y(Tag1[109]) );
  CLKINVX1 U561 ( .A(n578), .Y(Tag1[108]) );
  CLKINVX1 U562 ( .A(n579), .Y(Tag1[105]) );
  CLKINVX1 U563 ( .A(n580), .Y(Tag1[104]) );
  CLKINVX1 U564 ( .A(n581), .Y(Tag1[102]) );
  CLKINVX1 U565 ( .A(n582), .Y(Tag1[101]) );
  CLKINVX1 U566 ( .A(n583), .Y(Tag1[100]) );
  MXI2X1 U567 ( .A(n584), .B(n585), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_127_), .Y(n8213) );
  AOI21X1 U568 ( .A0(n586), .A1(n48), .B0(n70), .Y(n585) );
  CLKNAND2X2 U569 ( .A(n14), .B(n589), .Y(n584) );
  MXI2X1 U570 ( .A(n590), .B(n591), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_126_), .Y(n8212) );
  AOI21X1 U571 ( .A0(n592), .A1(n41), .B0(n75), .Y(n591) );
  NAND2BX1 U572 ( .AN(n592), .B(n33), .Y(n590) );
  MXI2X1 U573 ( .A(n593), .B(n594), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_125_), .Y(n8211) );
  AOI21X1 U574 ( .A0(n595), .A1(n41), .B0(n76), .Y(n594) );
  NAND2BX1 U575 ( .AN(n595), .B(n33), .Y(n593) );
  MXI2X1 U576 ( .A(n596), .B(n597), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_124_), .Y(n8210) );
  AOI21X1 U577 ( .A0(n598), .A1(n40), .B0(n76), .Y(n597) );
  NAND2BX1 U578 ( .AN(n598), .B(n34), .Y(n596) );
  MXI2X1 U579 ( .A(n599), .B(n600), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_123_), .Y(n8209) );
  AOI21X1 U580 ( .A0(n601), .A1(n40), .B0(n77), .Y(n600) );
  NAND2BX1 U581 ( .AN(n601), .B(n33), .Y(n599) );
  MXI2X1 U582 ( .A(n602), .B(n603), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_122_), .Y(n8208) );
  AOI21X1 U583 ( .A0(n604), .A1(n40), .B0(n77), .Y(n603) );
  NAND2BX1 U584 ( .AN(n604), .B(n34), .Y(n602) );
  MXI2X1 U585 ( .A(n605), .B(n606), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_121_), .Y(n8207) );
  AOI21X1 U586 ( .A0(n607), .A1(n40), .B0(n78), .Y(n606) );
  NAND2BX1 U587 ( .AN(n607), .B(n34), .Y(n605) );
  MXI2X1 U588 ( .A(n608), .B(n609), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_120_), .Y(n8206) );
  AOI21X1 U589 ( .A0(n610), .A1(n40), .B0(n79), .Y(n609) );
  NAND2BX1 U590 ( .AN(n610), .B(n34), .Y(n608) );
  MXI2X1 U591 ( .A(n611), .B(n612), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_119_), .Y(n8205) );
  AOI2B1X1 U592 ( .A1N(n613), .A0(n32), .B0(n82), .Y(n612) );
  CLKNAND2X2 U593 ( .A(n23), .B(n613), .Y(n611) );
  MXI2X1 U594 ( .A(n614), .B(n615), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_118_), .Y(n8204) );
  AOI21X1 U595 ( .A0(n616), .A1(n40), .B0(n80), .Y(n615) );
  CLKNAND2X2 U596 ( .A(n23), .B(n617), .Y(n614) );
  MXI2X1 U597 ( .A(n618), .B(n619), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_117_), .Y(n8203) );
  AOI21X1 U598 ( .A0(n620), .A1(n40), .B0(n80), .Y(n619) );
  CLKNAND2X2 U599 ( .A(n23), .B(n621), .Y(n618) );
  MXI2X1 U600 ( .A(n622), .B(n623), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_116_), .Y(n8202) );
  AOI21X1 U601 ( .A0(n624), .A1(n40), .B0(n81), .Y(n623) );
  CLKNAND2X2 U602 ( .A(n23), .B(n625), .Y(n622) );
  MXI2X1 U603 ( .A(n626), .B(n627), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_115_), .Y(n8201) );
  AOI21X1 U604 ( .A0(n628), .A1(n40), .B0(n82), .Y(n627) );
  CLKNAND2X2 U605 ( .A(n23), .B(n629), .Y(n626) );
  MXI2X1 U606 ( .A(n630), .B(n631), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_114_), .Y(n8200) );
  AOI21X1 U607 ( .A0(n632), .A1(n40), .B0(n65), .Y(n631) );
  CLKNAND2X2 U608 ( .A(n23), .B(n633), .Y(n630) );
  MXI2X1 U609 ( .A(n634), .B(n635), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_113_), .Y(n8199) );
  AOI21X1 U610 ( .A0(n636), .A1(n40), .B0(n66), .Y(n635) );
  CLKNAND2X2 U611 ( .A(n23), .B(n637), .Y(n634) );
  MXI2X1 U612 ( .A(n638), .B(n639), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_112_), .Y(n8198) );
  AOI21X1 U613 ( .A0(n640), .A1(n40), .B0(n67), .Y(n639) );
  CLKNAND2X2 U614 ( .A(n23), .B(n641), .Y(n638) );
  MXI2X1 U615 ( .A(n642), .B(n643), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_111_), .Y(n8197) );
  AOI2B1X1 U616 ( .A1N(n644), .A0(n32), .B0(n82), .Y(n643) );
  CLKNAND2X2 U617 ( .A(n23), .B(n644), .Y(n642) );
  MXI2X1 U618 ( .A(n645), .B(n646), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_110_), .Y(n8196) );
  AOI21X1 U619 ( .A0(n647), .A1(n39), .B0(n68), .Y(n646) );
  CLKNAND2X2 U620 ( .A(n23), .B(n648), .Y(n645) );
  MXI2X1 U621 ( .A(n649), .B(n650), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_109_), .Y(n8195) );
  AOI21X1 U622 ( .A0(n651), .A1(n39), .B0(n69), .Y(n650) );
  CLKNAND2X2 U623 ( .A(n23), .B(n652), .Y(n649) );
  MXI2X1 U624 ( .A(n653), .B(n654), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_108_), .Y(n8194) );
  AOI21X1 U625 ( .A0(n655), .A1(n39), .B0(n69), .Y(n654) );
  CLKNAND2X2 U626 ( .A(n24), .B(n656), .Y(n653) );
  MXI2X1 U627 ( .A(n657), .B(n658), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_107_), .Y(n8193) );
  AOI21X1 U628 ( .A0(n659), .A1(n39), .B0(n70), .Y(n658) );
  CLKNAND2X2 U629 ( .A(n24), .B(n660), .Y(n657) );
  MXI2X1 U630 ( .A(n661), .B(n662), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_106_), .Y(n8192) );
  AOI21X1 U631 ( .A0(n663), .A1(n39), .B0(n71), .Y(n662) );
  CLKNAND2X2 U632 ( .A(n24), .B(n664), .Y(n661) );
  MXI2X1 U633 ( .A(n665), .B(n666), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_105_), .Y(n8191) );
  AOI21X1 U634 ( .A0(n667), .A1(n39), .B0(n72), .Y(n666) );
  CLKNAND2X2 U635 ( .A(n24), .B(n668), .Y(n665) );
  MXI2X1 U636 ( .A(n669), .B(n670), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_104_), .Y(n8190) );
  AOI21X1 U637 ( .A0(n671), .A1(n39), .B0(n72), .Y(n670) );
  CLKNAND2X2 U638 ( .A(n24), .B(n672), .Y(n669) );
  MXI2X1 U639 ( .A(n673), .B(n674), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_103_), .Y(n8189) );
  AOI2B1X1 U640 ( .A1N(n675), .A0(n31), .B0(n82), .Y(n674) );
  CLKNAND2X2 U641 ( .A(n24), .B(n675), .Y(n673) );
  MXI2X1 U642 ( .A(n676), .B(n677), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_102_), .Y(n8188) );
  AOI21X1 U643 ( .A0(n678), .A1(n39), .B0(n73), .Y(n677) );
  CLKNAND2X2 U644 ( .A(n27), .B(n679), .Y(n676) );
  MXI2X1 U645 ( .A(n680), .B(n681), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_101_), .Y(n8187) );
  AOI21X1 U646 ( .A0(n682), .A1(n38), .B0(n65), .Y(n681) );
  CLKNAND2X2 U647 ( .A(n25), .B(n683), .Y(n680) );
  MXI2X1 U648 ( .A(n684), .B(n685), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_100_), .Y(n8186) );
  AOI21X1 U649 ( .A0(n686), .A1(n38), .B0(n73), .Y(n685) );
  CLKNAND2X2 U650 ( .A(n25), .B(n687), .Y(n684) );
  MXI2X1 U651 ( .A(n688), .B(n689), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_99_), .Y(n8185) );
  AOI21X1 U652 ( .A0(n690), .A1(n38), .B0(n73), .Y(n689) );
  CLKNAND2X2 U653 ( .A(n25), .B(n691), .Y(n688) );
  MXI2X1 U654 ( .A(n692), .B(n693), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_98_), .Y(n8184) );
  AOI21X1 U655 ( .A0(n694), .A1(n38), .B0(n73), .Y(n693) );
  CLKNAND2X2 U656 ( .A(n25), .B(n695), .Y(n692) );
  MXI2X1 U657 ( .A(n696), .B(n697), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_97_), .Y(n8183) );
  AOI21X1 U658 ( .A0(n698), .A1(n38), .B0(n73), .Y(n697) );
  CLKNAND2X2 U659 ( .A(n25), .B(n699), .Y(n696) );
  MXI2X1 U660 ( .A(n700), .B(n701), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_96_), .Y(n8182) );
  AOI21X1 U661 ( .A0(n702), .A1(n38), .B0(n73), .Y(n701) );
  CLKNAND2X2 U662 ( .A(n25), .B(n703), .Y(n700) );
  MXI2X1 U663 ( .A(n704), .B(n705), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_95_), .Y(n8181) );
  AOI2B1X1 U664 ( .A1N(n706), .A0(n32), .B0(n82), .Y(n705) );
  CLKNAND2X2 U665 ( .A(n26), .B(n706), .Y(n704) );
  MXI2X1 U666 ( .A(n707), .B(n708), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_94_), .Y(n8180) );
  AOI21X1 U667 ( .A0(n709), .A1(n38), .B0(n73), .Y(n708) );
  CLKNAND2X2 U668 ( .A(n26), .B(n710), .Y(n707) );
  MXI2X1 U669 ( .A(n711), .B(n712), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_93_), .Y(n8179) );
  AOI21X1 U670 ( .A0(n713), .A1(n38), .B0(n73), .Y(n712) );
  CLKNAND2X2 U671 ( .A(n26), .B(n714), .Y(n711) );
  MXI2X1 U672 ( .A(n715), .B(n716), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_92_), .Y(n8178) );
  AOI21X1 U673 ( .A0(n717), .A1(n37), .B0(n73), .Y(n716) );
  CLKNAND2X2 U674 ( .A(n26), .B(n718), .Y(n715) );
  MXI2X1 U675 ( .A(n719), .B(n720), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_91_), .Y(n8177) );
  AOI21X1 U676 ( .A0(n721), .A1(n37), .B0(n73), .Y(n720) );
  CLKNAND2X2 U677 ( .A(n26), .B(n722), .Y(n719) );
  MXI2X1 U678 ( .A(n723), .B(n724), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_90_), .Y(n8176) );
  AOI21X1 U679 ( .A0(n725), .A1(n37), .B0(n73), .Y(n724) );
  CLKNAND2X2 U680 ( .A(n26), .B(n726), .Y(n723) );
  MXI2X1 U681 ( .A(n727), .B(n728), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_89_), .Y(n8175) );
  AOI21X1 U682 ( .A0(n729), .A1(n37), .B0(n72), .Y(n728) );
  CLKNAND2X2 U683 ( .A(n27), .B(n730), .Y(n727) );
  MXI2X1 U684 ( .A(n731), .B(n732), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_88_), .Y(n8174) );
  AOI21X1 U685 ( .A0(n733), .A1(n37), .B0(n72), .Y(n732) );
  CLKNAND2X2 U686 ( .A(n27), .B(n734), .Y(n731) );
  MXI2X1 U687 ( .A(n735), .B(n736), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_87_), .Y(n8173) );
  AOI2B1X1 U688 ( .A1N(n737), .A0(n31), .B0(n83), .Y(n736) );
  CLKNAND2X2 U689 ( .A(n27), .B(n737), .Y(n735) );
  MXI2X1 U690 ( .A(n738), .B(n739), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_86_), .Y(n8172) );
  AOI21X1 U691 ( .A0(n740), .A1(n37), .B0(n72), .Y(n739) );
  CLKNAND2X2 U692 ( .A(n27), .B(n741), .Y(n738) );
  MXI2X1 U693 ( .A(n742), .B(n743), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_85_), .Y(n8171) );
  AOI21X1 U694 ( .A0(n744), .A1(n37), .B0(n72), .Y(n743) );
  CLKNAND2X2 U695 ( .A(n27), .B(n745), .Y(n742) );
  MXI2X1 U696 ( .A(n746), .B(n747), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_84_), .Y(n8170) );
  AOI21X1 U697 ( .A0(n748), .A1(n36), .B0(n72), .Y(n747) );
  CLKNAND2X2 U698 ( .A(n28), .B(n749), .Y(n746) );
  MXI2X1 U699 ( .A(n750), .B(n751), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_83_), .Y(n8169) );
  AOI21X1 U700 ( .A0(n752), .A1(n37), .B0(n72), .Y(n751) );
  CLKNAND2X2 U701 ( .A(n28), .B(n753), .Y(n750) );
  MXI2X1 U702 ( .A(n754), .B(n755), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_82_), .Y(n8168) );
  AOI21X1 U703 ( .A0(n756), .A1(n36), .B0(n72), .Y(n755) );
  CLKNAND2X2 U704 ( .A(n28), .B(n757), .Y(n754) );
  MXI2X1 U705 ( .A(n758), .B(n759), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_81_), .Y(n8167) );
  AOI21X1 U706 ( .A0(n760), .A1(n36), .B0(n72), .Y(n759) );
  CLKNAND2X2 U707 ( .A(n28), .B(n761), .Y(n758) );
  MXI2X1 U708 ( .A(n762), .B(n763), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_80_), .Y(n8166) );
  AOI21X1 U709 ( .A0(n764), .A1(n36), .B0(n72), .Y(n763) );
  CLKNAND2X2 U710 ( .A(n28), .B(n765), .Y(n762) );
  MXI2X1 U711 ( .A(n766), .B(n767), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_79_), .Y(n8165) );
  AOI2B1X1 U712 ( .A1N(n768), .A0(n31), .B0(n83), .Y(n767) );
  CLKNAND2X2 U713 ( .A(n28), .B(n768), .Y(n766) );
  MXI2X1 U714 ( .A(n769), .B(n770), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_78_), .Y(n8164) );
  AOI21X1 U715 ( .A0(n771), .A1(n36), .B0(n72), .Y(n770) );
  CLKNAND2X2 U716 ( .A(n28), .B(n772), .Y(n769) );
  MXI2X1 U717 ( .A(n773), .B(n774), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_77_), .Y(n8163) );
  AOI21X1 U718 ( .A0(n775), .A1(n36), .B0(n72), .Y(n774) );
  CLKNAND2X2 U719 ( .A(n28), .B(n776), .Y(n773) );
  MXI2X1 U720 ( .A(n777), .B(n778), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_76_), .Y(n8162) );
  AOI21X1 U721 ( .A0(n779), .A1(n36), .B0(n71), .Y(n778) );
  CLKNAND2X2 U722 ( .A(n29), .B(n780), .Y(n777) );
  MXI2X1 U723 ( .A(n781), .B(n782), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_75_), .Y(n8161) );
  AOI21X1 U724 ( .A0(n783), .A1(n35), .B0(n71), .Y(n782) );
  CLKNAND2X2 U725 ( .A(n29), .B(n784), .Y(n781) );
  MXI2X1 U726 ( .A(n785), .B(n786), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_74_), .Y(n8160) );
  AOI21X1 U727 ( .A0(n787), .A1(n35), .B0(n71), .Y(n786) );
  CLKNAND2X2 U728 ( .A(n29), .B(n788), .Y(n785) );
  MXI2X1 U729 ( .A(n789), .B(n790), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_73_), .Y(n8159) );
  AOI21X1 U730 ( .A0(n791), .A1(n35), .B0(n71), .Y(n790) );
  CLKNAND2X2 U731 ( .A(n30), .B(n792), .Y(n789) );
  MXI2X1 U732 ( .A(n793), .B(n794), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_72_), .Y(n8158) );
  AOI21X1 U733 ( .A0(n795), .A1(n35), .B0(n71), .Y(n794) );
  CLKNAND2X2 U734 ( .A(n30), .B(n796), .Y(n793) );
  MXI2X1 U735 ( .A(n797), .B(n798), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_71_), .Y(n8157) );
  AOI2B1X1 U736 ( .A1N(n799), .A0(n32), .B0(n83), .Y(n798) );
  CLKNAND2X2 U737 ( .A(n29), .B(n799), .Y(n797) );
  MXI2X1 U738 ( .A(n800), .B(n801), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_70_), .Y(n8156) );
  AOI21X1 U739 ( .A0(n802), .A1(n35), .B0(n71), .Y(n801) );
  CLKNAND2X2 U740 ( .A(n30), .B(n803), .Y(n800) );
  MXI2X1 U741 ( .A(n804), .B(n805), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_69_), .Y(n8155) );
  AOI21X1 U742 ( .A0(n806), .A1(n35), .B0(n71), .Y(n805) );
  CLKNAND2X2 U743 ( .A(n31), .B(n807), .Y(n804) );
  MXI2X1 U744 ( .A(n808), .B(n809), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_68_), .Y(n8154) );
  AOI21X1 U745 ( .A0(n810), .A1(n35), .B0(n71), .Y(n809) );
  CLKNAND2X2 U746 ( .A(n30), .B(n811), .Y(n808) );
  MXI2X1 U747 ( .A(n812), .B(n813), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_67_), .Y(n8153) );
  AOI21X1 U748 ( .A0(n814), .A1(n35), .B0(n71), .Y(n813) );
  CLKNAND2X2 U749 ( .A(n30), .B(n815), .Y(n812) );
  MXI2X1 U750 ( .A(n816), .B(n817), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_66_), .Y(n8152) );
  AOI21X1 U751 ( .A0(n818), .A1(n48), .B0(n71), .Y(n817) );
  CLKNAND2X2 U752 ( .A(n31), .B(n819), .Y(n816) );
  MXI2X1 U753 ( .A(n820), .B(n821), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_65_), .Y(n8151) );
  AOI21X1 U754 ( .A0(n822), .A1(n48), .B0(n71), .Y(n821) );
  CLKNAND2X2 U755 ( .A(n31), .B(n823), .Y(n820) );
  MXI2X1 U756 ( .A(n824), .B(n825), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_64_), .Y(n8150) );
  AOI21X1 U757 ( .A0(n826), .A1(n48), .B0(n71), .Y(n825) );
  CLKNAND2X2 U758 ( .A(n30), .B(n827), .Y(n824) );
  MXI2X1 U759 ( .A(n828), .B(n829), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_63_), .Y(n8149) );
  AOI2B1X1 U760 ( .A1N(n830), .A0(n32), .B0(n82), .Y(n829) );
  CLKNAND2X2 U761 ( .A(n31), .B(n830), .Y(n828) );
  MXI2X1 U762 ( .A(n831), .B(n832), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_62_), .Y(n8148) );
  AOI21X1 U763 ( .A0(n833), .A1(n47), .B0(n70), .Y(n832) );
  CLKNAND2X2 U764 ( .A(n29), .B(n834), .Y(n831) );
  MXI2X1 U765 ( .A(n835), .B(n836), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_61_), .Y(n8147) );
  AOI21X1 U766 ( .A0(n837), .A1(n47), .B0(n70), .Y(n836) );
  CLKNAND2X2 U767 ( .A(n14), .B(n838), .Y(n835) );
  MXI2X1 U768 ( .A(n839), .B(n840), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_60_), .Y(n8146) );
  AOI21X1 U769 ( .A0(n841), .A1(n47), .B0(n70), .Y(n840) );
  CLKNAND2X2 U770 ( .A(n14), .B(n842), .Y(n839) );
  MXI2X1 U771 ( .A(n843), .B(n844), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_59_), .Y(n8145) );
  AOI21X1 U772 ( .A0(n845), .A1(n47), .B0(n70), .Y(n844) );
  CLKNAND2X2 U773 ( .A(n14), .B(n846), .Y(n843) );
  MXI2X1 U774 ( .A(n847), .B(n848), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_58_), .Y(n8144) );
  AOI21X1 U775 ( .A0(n849), .A1(n47), .B0(n70), .Y(n848) );
  CLKNAND2X2 U776 ( .A(n14), .B(n850), .Y(n847) );
  MXI2X1 U777 ( .A(n851), .B(n852), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_57_), .Y(n8143) );
  AOI21X1 U778 ( .A0(n853), .A1(n47), .B0(n70), .Y(n852) );
  CLKNAND2X2 U779 ( .A(n14), .B(n854), .Y(n851) );
  MXI2X1 U780 ( .A(n855), .B(n856), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_56_), .Y(n8142) );
  AOI21X1 U781 ( .A0(n857), .A1(n47), .B0(n70), .Y(n856) );
  CLKNAND2X2 U782 ( .A(n14), .B(n858), .Y(n855) );
  MXI2X1 U783 ( .A(n859), .B(n860), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_55_), .Y(n8141) );
  AOI2B1X1 U784 ( .A1N(n861), .A0(n32), .B0(n83), .Y(n860) );
  CLKNAND2X2 U785 ( .A(n15), .B(n861), .Y(n859) );
  MXI2X1 U786 ( .A(n862), .B(n863), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_54_), .Y(n8140) );
  AOI21X1 U787 ( .A0(n864), .A1(n47), .B0(n70), .Y(n863) );
  CLKNAND2X2 U788 ( .A(n15), .B(n865), .Y(n862) );
  MXI2X1 U789 ( .A(n866), .B(n867), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_53_), .Y(n8139) );
  AOI21X1 U790 ( .A0(n868), .A1(n46), .B0(n70), .Y(n867) );
  CLKNAND2X2 U791 ( .A(n15), .B(n869), .Y(n866) );
  MXI2X1 U792 ( .A(n870), .B(n871), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_52_), .Y(n8138) );
  AOI21X1 U793 ( .A0(n872), .A1(n46), .B0(n70), .Y(n871) );
  CLKNAND2X2 U794 ( .A(n15), .B(n873), .Y(n870) );
  MXI2X1 U795 ( .A(n874), .B(n875), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_51_), .Y(n8137) );
  AOI21X1 U796 ( .A0(n876), .A1(n46), .B0(n70), .Y(n875) );
  CLKNAND2X2 U797 ( .A(n15), .B(n877), .Y(n874) );
  MXI2X1 U798 ( .A(n878), .B(n879), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_50_), .Y(n8136) );
  AOI21X1 U799 ( .A0(n880), .A1(n46), .B0(n69), .Y(n879) );
  CLKNAND2X2 U800 ( .A(n15), .B(n881), .Y(n878) );
  MXI2X1 U801 ( .A(n882), .B(n883), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_49_), .Y(n8135) );
  AOI21X1 U802 ( .A0(n884), .A1(n46), .B0(n69), .Y(n883) );
  CLKNAND2X2 U803 ( .A(n16), .B(n885), .Y(n882) );
  MXI2X1 U804 ( .A(n886), .B(n887), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_48_), .Y(n8134) );
  AOI21X1 U805 ( .A0(n888), .A1(n46), .B0(n69), .Y(n887) );
  CLKNAND2X2 U806 ( .A(n16), .B(n889), .Y(n886) );
  MXI2X1 U807 ( .A(n890), .B(n891), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_47_), .Y(n8133) );
  AOI2B1X1 U808 ( .A1N(n892), .A0(n32), .B0(n83), .Y(n891) );
  CLKNAND2X2 U809 ( .A(n16), .B(n892), .Y(n890) );
  MXI2X1 U810 ( .A(n893), .B(n894), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_46_), .Y(n8132) );
  AOI21X1 U811 ( .A0(n895), .A1(n46), .B0(n69), .Y(n894) );
  CLKNAND2X2 U812 ( .A(n16), .B(n896), .Y(n893) );
  MXI2X1 U813 ( .A(n897), .B(n898), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_45_), .Y(n8131) );
  AOI21X1 U814 ( .A0(n899), .A1(n46), .B0(n69), .Y(n898) );
  CLKNAND2X2 U815 ( .A(n16), .B(n900), .Y(n897) );
  MXI2X1 U816 ( .A(n901), .B(n902), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_44_), .Y(n8130) );
  AOI21X1 U817 ( .A0(n903), .A1(n45), .B0(n69), .Y(n902) );
  CLKNAND2X2 U818 ( .A(n16), .B(n904), .Y(n901) );
  MXI2X1 U819 ( .A(n905), .B(n906), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_43_), .Y(n8129) );
  AOI21X1 U820 ( .A0(n907), .A1(n45), .B0(n69), .Y(n906) );
  CLKNAND2X2 U821 ( .A(n17), .B(n908), .Y(n905) );
  MXI2X1 U822 ( .A(n909), .B(n910), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_42_), .Y(n8128) );
  AOI21X1 U823 ( .A0(n911), .A1(n45), .B0(n69), .Y(n910) );
  CLKNAND2X2 U824 ( .A(n17), .B(n912), .Y(n909) );
  MXI2X1 U825 ( .A(n913), .B(n914), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_41_), .Y(n8127) );
  AOI21X1 U826 ( .A0(n915), .A1(n45), .B0(n69), .Y(n914) );
  CLKNAND2X2 U827 ( .A(n17), .B(n916), .Y(n913) );
  MXI2X1 U828 ( .A(n917), .B(n918), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_40_), .Y(n8126) );
  AOI21X1 U829 ( .A0(n919), .A1(n45), .B0(n69), .Y(n918) );
  CLKNAND2X2 U830 ( .A(n17), .B(n920), .Y(n917) );
  MXI2X1 U831 ( .A(n921), .B(n922), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_39_), .Y(n8125) );
  AOI2B1X1 U832 ( .A1N(n923), .A0(n31), .B0(n83), .Y(n922) );
  CLKNAND2X2 U833 ( .A(n17), .B(n923), .Y(n921) );
  MXI2X1 U834 ( .A(n924), .B(n925), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_38_), .Y(n8124) );
  AOI21X1 U835 ( .A0(n926), .A1(n45), .B0(n68), .Y(n925) );
  CLKNAND2X2 U836 ( .A(n17), .B(n927), .Y(n924) );
  MXI2X1 U837 ( .A(n928), .B(n929), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_37_), .Y(n8123) );
  AOI21X1 U838 ( .A0(n930), .A1(n45), .B0(n68), .Y(n929) );
  CLKNAND2X2 U839 ( .A(n18), .B(n931), .Y(n928) );
  MXI2X1 U840 ( .A(n932), .B(n933), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_36_), .Y(n8122) );
  AOI21X1 U841 ( .A0(n934), .A1(n45), .B0(n68), .Y(n933) );
  CLKNAND2X2 U842 ( .A(n18), .B(n935), .Y(n932) );
  MXI2X1 U843 ( .A(n936), .B(n937), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_35_), .Y(n8121) );
  AOI21X1 U844 ( .A0(n938), .A1(n45), .B0(n68), .Y(n937) );
  CLKNAND2X2 U845 ( .A(n18), .B(n939), .Y(n936) );
  MXI2X1 U846 ( .A(n940), .B(n941), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_34_), .Y(n8120) );
  AOI21X1 U847 ( .A0(n942), .A1(n44), .B0(n68), .Y(n941) );
  CLKNAND2X2 U848 ( .A(n18), .B(n943), .Y(n940) );
  MXI2X1 U849 ( .A(n944), .B(n945), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_33_), .Y(n8119) );
  AOI21X1 U850 ( .A0(n946), .A1(n44), .B0(n68), .Y(n945) );
  CLKNAND2X2 U851 ( .A(n18), .B(n947), .Y(n944) );
  MXI2X1 U852 ( .A(n948), .B(n949), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_32_), .Y(n8118) );
  AOI21X1 U853 ( .A0(n950), .A1(n44), .B0(n68), .Y(n949) );
  CLKNAND2X2 U854 ( .A(n18), .B(n951), .Y(n948) );
  MXI2X1 U855 ( .A(n952), .B(n953), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_31_), .Y(n8117) );
  AOI2B1X1 U856 ( .A1N(n954), .A0(n31), .B0(n83), .Y(n953) );
  CLKNAND2X2 U857 ( .A(n19), .B(n954), .Y(n952) );
  MXI2X1 U858 ( .A(n955), .B(n956), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_30_), .Y(n8116) );
  AOI21X1 U859 ( .A0(n957), .A1(n44), .B0(n68), .Y(n956) );
  CLKNAND2X2 U860 ( .A(n19), .B(n958), .Y(n955) );
  MXI2X1 U861 ( .A(n959), .B(n960), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_29_), .Y(n8115) );
  AOI21X1 U862 ( .A0(n961), .A1(n44), .B0(n68), .Y(n960) );
  CLKNAND2X2 U863 ( .A(n19), .B(n962), .Y(n959) );
  MXI2X1 U864 ( .A(n963), .B(n964), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_28_), .Y(n8114) );
  AOI21X1 U865 ( .A0(n965), .A1(n44), .B0(n68), .Y(n964) );
  CLKNAND2X2 U866 ( .A(n19), .B(n966), .Y(n963) );
  MXI2X1 U867 ( .A(n967), .B(n968), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_27_), .Y(n8113) );
  AOI21X1 U868 ( .A0(n969), .A1(n44), .B0(n68), .Y(n968) );
  CLKNAND2X2 U869 ( .A(n19), .B(n970), .Y(n967) );
  MXI2X1 U870 ( .A(n971), .B(n972), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_26_), .Y(n8112) );
  AOI21X1 U871 ( .A0(n973), .A1(n43), .B0(n68), .Y(n972) );
  CLKNAND2X2 U872 ( .A(n19), .B(n974), .Y(n971) );
  MXI2X1 U873 ( .A(n975), .B(n976), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_25_), .Y(n8111) );
  AOI21X1 U874 ( .A0(n977), .A1(n43), .B0(n67), .Y(n976) );
  CLKNAND2X2 U875 ( .A(n20), .B(n978), .Y(n975) );
  MXI2X1 U876 ( .A(n979), .B(n980), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_24_), .Y(n8110) );
  AOI21X1 U877 ( .A0(n981), .A1(n43), .B0(n67), .Y(n980) );
  CLKNAND2X2 U878 ( .A(n20), .B(n982), .Y(n979) );
  MXI2X1 U879 ( .A(n983), .B(n984), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_23_), .Y(n8109) );
  AOI2B1X1 U880 ( .A1N(n985), .A0(n31), .B0(n83), .Y(n984) );
  CLKNAND2X2 U881 ( .A(n20), .B(n985), .Y(n983) );
  MXI2X1 U882 ( .A(n986), .B(n987), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_22_), .Y(n8108) );
  AOI21X1 U883 ( .A0(n988), .A1(n43), .B0(n67), .Y(n987) );
  CLKNAND2X2 U884 ( .A(n20), .B(n989), .Y(n986) );
  MXI2X1 U885 ( .A(n990), .B(n991), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_21_), .Y(n8107) );
  AOI21X1 U886 ( .A0(n992), .A1(n43), .B0(n67), .Y(n991) );
  CLKNAND2X2 U887 ( .A(n20), .B(n993), .Y(n990) );
  MXI2X1 U888 ( .A(n994), .B(n995), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_20_), .Y(n8106) );
  AOI21X1 U889 ( .A0(n996), .A1(n43), .B0(n67), .Y(n995) );
  CLKNAND2X2 U890 ( .A(n20), .B(n997), .Y(n994) );
  MXI2X1 U891 ( .A(n998), .B(n999), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_19_), .Y(n8105) );
  AOI21X1 U892 ( .A0(n1000), .A1(n43), .B0(n67), .Y(n999) );
  CLKNAND2X2 U893 ( .A(n21), .B(n1001), .Y(n998) );
  MXI2X1 U894 ( .A(n1002), .B(n1003), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_18_), .Y(n8104) );
  AOI21X1 U895 ( .A0(n1004), .A1(n43), .B0(n67), .Y(n1003) );
  CLKNAND2X2 U896 ( .A(n21), .B(n1005), .Y(n1002) );
  MXI2X1 U897 ( .A(n1006), .B(n1007), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_17_), .Y(n8103) );
  AOI21X1 U898 ( .A0(n1008), .A1(n43), .B0(n67), .Y(n1007) );
  CLKNAND2X2 U899 ( .A(n21), .B(n1009), .Y(n1006) );
  MXI2X1 U900 ( .A(n1010), .B(n1011), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_16_), .Y(n8102) );
  AOI21X1 U901 ( .A0(n1012), .A1(n42), .B0(n67), .Y(n1011) );
  CLKNAND2X2 U902 ( .A(n21), .B(n1013), .Y(n1010) );
  MXI2X1 U903 ( .A(n1014), .B(n1015), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_15_), .Y(n8101) );
  AOI2B1X1 U904 ( .A1N(n1016), .A0(n31), .B0(n83), .Y(n1015) );
  CLKNAND2X2 U905 ( .A(n21), .B(n1016), .Y(n1014) );
  MXI2X1 U906 ( .A(n1017), .B(n1018), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_14_), .Y(n8100) );
  AOI21X1 U907 ( .A0(n1019), .A1(n42), .B0(n67), .Y(n1018) );
  CLKNAND2X2 U908 ( .A(n21), .B(n1020), .Y(n1017) );
  MXI2X1 U909 ( .A(n1021), .B(n1022), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_13_), .Y(n8099) );
  AOI21X1 U910 ( .A0(n1023), .A1(n42), .B0(n67), .Y(n1022) );
  CLKNAND2X2 U911 ( .A(n22), .B(n1024), .Y(n1021) );
  MXI2X1 U912 ( .A(n1025), .B(n1026), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_12_), .Y(n8098) );
  AOI21X1 U913 ( .A0(n1027), .A1(n42), .B0(n67), .Y(n1026) );
  CLKNAND2X2 U914 ( .A(n22), .B(n1028), .Y(n1025) );
  MXI2X1 U915 ( .A(n1029), .B(n1030), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_11_), .Y(n8097) );
  AOI21X1 U916 ( .A0(n1031), .A1(n42), .B0(n66), .Y(n1030) );
  CLKNAND2X2 U917 ( .A(n22), .B(n1032), .Y(n1029) );
  MXI2X1 U918 ( .A(n1033), .B(n1034), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_10_), .Y(n8096) );
  AOI21X1 U919 ( .A0(n1035), .A1(n42), .B0(n66), .Y(n1034) );
  CLKNAND2X2 U920 ( .A(n22), .B(n1036), .Y(n1033) );
  MXI2X1 U921 ( .A(n1037), .B(n1038), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_9_), .Y(n8095) );
  AOI21X1 U922 ( .A0(n1039), .A1(n42), .B0(n66), .Y(n1038) );
  CLKNAND2X2 U923 ( .A(n22), .B(n1040), .Y(n1037) );
  MXI2X1 U924 ( .A(n1041), .B(n1042), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_8_), .Y(n8094) );
  AOI21X1 U925 ( .A0(n1043), .A1(n42), .B0(n66), .Y(n1042) );
  CLKNAND2X2 U926 ( .A(n22), .B(n1044), .Y(n1041) );
  MXI2X1 U927 ( .A(n1045), .B(n1046), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_7_), .Y(n8093) );
  AOI2B1X1 U928 ( .A1N(n1047), .A0(n32), .B0(n83), .Y(n1046) );
  CLKNAND2X2 U929 ( .A(n22), .B(n1047), .Y(n1045) );
  MXI2X1 U930 ( .A(n1048), .B(n1049), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_6_), .Y(n8092) );
  AOI21X1 U931 ( .A0(n1050), .A1(n41), .B0(n66), .Y(n1049) );
  NAND2BX1 U932 ( .AN(n1050), .B(n34), .Y(n1048) );
  MXI2X1 U933 ( .A(n1051), .B(n1052), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_5_), .Y(n8091) );
  AOI21X1 U934 ( .A0(n1053), .A1(n41), .B0(n66), .Y(n1052) );
  NAND2BX1 U935 ( .AN(n1053), .B(n34), .Y(n1051) );
  MXI2X1 U936 ( .A(n1054), .B(n1055), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_4_), .Y(n8090) );
  AOI21X1 U937 ( .A0(n1056), .A1(n41), .B0(n66), .Y(n1055) );
  NAND2BX1 U938 ( .AN(n1056), .B(n34), .Y(n1054) );
  MXI2X1 U939 ( .A(n1057), .B(n1058), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_3_), .Y(n8089) );
  AOI21X1 U940 ( .A0(n1059), .A1(n41), .B0(n66), .Y(n1058) );
  NAND2BX1 U941 ( .AN(n1059), .B(n33), .Y(n1057) );
  MXI2X1 U942 ( .A(n1060), .B(n1061), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_2_), .Y(n8088) );
  AOI21X1 U943 ( .A0(n1062), .A1(n41), .B0(n66), .Y(n1061) );
  NAND2BX1 U944 ( .AN(n1062), .B(n34), .Y(n1060) );
  MXI2X1 U945 ( .A(n1063), .B(n1064), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_1_), .Y(n8087) );
  AOI21X1 U946 ( .A0(n1065), .A1(n41), .B0(n66), .Y(n1064) );
  NAND2BX1 U947 ( .AN(n1065), .B(n33), .Y(n1063) );
  MXI2X1 U948 ( .A(n1066), .B(n1067), .S0(
        Inst_forkAE_MainPart2_Tag_Reg_Output_0_), .Y(n8086) );
  AOI21X1 U949 ( .A0(n1068), .A1(n41), .B0(n66), .Y(n1067) );
  NAND2BX1 U950 ( .AN(n1068), .B(n33), .Y(n1066) );
  OAI2B2X1 U951 ( .A1N(Tag2[127]), .A0(n103), .B0(n1070), .B1(n132), .Y(n7829)
         );
  CLKINVX1 U952 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[127]), .Y(n1070) );
  XOR2X1 U953 ( .A(n1072), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[127]), .Y(
        Tag2[127]) );
  OAI2B2X1 U954 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[126]), .A0(n126), 
        .B0(n517), .B1(n108), .Y(n7828) );
  XOR2X1 U955 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[126]), .B(n1073), .Y(
        n517) );
  OAI2B2X1 U956 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[125]), .A0(n126), 
        .B0(n518), .B1(n108), .Y(n7827) );
  XOR2X1 U957 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[125]), .B(n1074), .Y(
        n518) );
  OAI2B2X1 U958 ( .A1N(Tag2[124]), .A0(n96), .B0(n1075), .B1(n132), .Y(n7826)
         );
  CLKINVX1 U959 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[124]), .Y(n1075) );
  XOR2X1 U960 ( .A(n1076), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[124]), .Y(
        Tag2[124]) );
  OAI2B2X1 U961 ( .A1N(Tag2[123]), .A0(n96), .B0(n1077), .B1(n132), .Y(n7825)
         );
  CLKINVX1 U962 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[123]), .Y(n1077) );
  XOR2X1 U963 ( .A(n1078), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[123]), .Y(
        Tag2[123]) );
  OAI2B2X1 U964 ( .A1N(Tag2[122]), .A0(n96), .B0(n1079), .B1(n131), .Y(n7824)
         );
  CLKINVX1 U965 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[122]), .Y(n1079) );
  XOR2X1 U966 ( .A(n1080), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[122]), .Y(
        Tag2[122]) );
  OAI2B2X1 U967 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[121]), .A0(n127), 
        .B0(n519), .B1(n109), .Y(n7823) );
  XOR2X1 U968 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[121]), .B(n1081), .Y(
        n519) );
  OAI2B2X1 U969 ( .A1N(Tag2[120]), .A0(n96), .B0(n1082), .B1(n131), .Y(n7822)
         );
  CLKINVX1 U970 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[120]), .Y(n1082) );
  XOR2X1 U971 ( .A(n1083), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[120]), .Y(
        Tag2[120]) );
  OAI2B2X1 U972 ( .A1N(Tag2[119]), .A0(n96), .B0(n1084), .B1(n131), .Y(n7821)
         );
  CLKINVX1 U973 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[119]), .Y(n1084) );
  XOR2X1 U974 ( .A(n1085), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[119]), .Y(
        Tag2[119]) );
  OAI2B2X1 U975 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[118]), .A0(n127), 
        .B0(n520), .B1(n108), .Y(n7820) );
  XOR2X1 U976 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[118]), .B(n1086), .Y(
        n520) );
  OAI2B2X1 U977 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[117]), .A0(n128), 
        .B0(n521), .B1(n109), .Y(n7819) );
  XOR2X1 U978 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[117]), .B(n1087), .Y(
        n521) );
  OAI2B2X1 U979 ( .A1N(Tag2[116]), .A0(n96), .B0(n1088), .B1(n131), .Y(n7818)
         );
  CLKINVX1 U980 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[116]), .Y(n1088) );
  XOR2X1 U981 ( .A(n1089), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[116]), .Y(
        Tag2[116]) );
  OAI2B2X1 U982 ( .A1N(Tag2[115]), .A0(n96), .B0(n1090), .B1(n131), .Y(n7817)
         );
  CLKINVX1 U983 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[115]), .Y(n1090) );
  XOR2X1 U984 ( .A(n1091), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[115]), .Y(
        Tag2[115]) );
  OAI2B2X1 U985 ( .A1N(Tag2[114]), .A0(n96), .B0(n1092), .B1(n131), .Y(n7816)
         );
  CLKINVX1 U986 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[114]), .Y(n1092) );
  XOR2X1 U987 ( .A(n1093), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[114]), .Y(
        Tag2[114]) );
  OAI2B2X1 U988 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[113]), .A0(n127), 
        .B0(n522), .B1(n108), .Y(n7815) );
  XOR2X1 U989 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[113]), .B(n1094), .Y(
        n522) );
  OAI2B2X1 U990 ( .A1N(Tag2[112]), .A0(n96), .B0(n1095), .B1(n130), .Y(n7814)
         );
  CLKINVX1 U991 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[112]), .Y(n1095) );
  XOR2X1 U992 ( .A(n1096), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[112]), .Y(
        Tag2[112]) );
  OAI2B2X1 U993 ( .A1N(Tag2[111]), .A0(n96), .B0(n1097), .B1(n130), .Y(n7813)
         );
  CLKINVX1 U994 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[111]), .Y(n1097) );
  XOR2X1 U995 ( .A(n1098), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[111]), .Y(
        Tag2[111]) );
  OAI2B2X1 U996 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[110]), .A0(n127), 
        .B0(n523), .B1(n109), .Y(n7812) );
  XOR2X1 U997 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[110]), .B(n1099), .Y(
        n523) );
  OAI2B2X1 U998 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[109]), .A0(n127), 
        .B0(n524), .B1(n109), .Y(n7811) );
  XOR2X1 U999 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[109]), .B(n1100), .Y(
        n524) );
  OAI2B2X1 U1000 ( .A1N(Tag2[108]), .A0(n96), .B0(n1101), .B1(n130), .Y(n7810)
         );
  CLKINVX1 U1001 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[108]), .Y(n1101)
         );
  XOR2X1 U1002 ( .A(n1102), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[108]), 
        .Y(Tag2[108]) );
  OAI2B2X1 U1003 ( .A1N(Tag2[107]), .A0(n96), .B0(n1103), .B1(n130), .Y(n7809)
         );
  CLKINVX1 U1004 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[107]), .Y(n1103)
         );
  XOR2X1 U1005 ( .A(n1104), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[107]), 
        .Y(Tag2[107]) );
  OAI2B2X1 U1006 ( .A1N(Tag2[106]), .A0(n97), .B0(n1105), .B1(n130), .Y(n7808)
         );
  CLKINVX1 U1007 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[106]), .Y(n1105)
         );
  XOR2X1 U1008 ( .A(n1106), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[106]), 
        .Y(Tag2[106]) );
  OAI2B2X1 U1009 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[105]), .A0(n127), 
        .B0(n525), .B1(n110), .Y(n7807) );
  XOR2X1 U1010 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[105]), .B(n1107), 
        .Y(n525) );
  OAI2B2X1 U1011 ( .A1N(Tag2[104]), .A0(n97), .B0(n1108), .B1(n130), .Y(n7806)
         );
  CLKINVX1 U1012 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[104]), .Y(n1108)
         );
  XOR2X1 U1013 ( .A(n1109), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[104]), 
        .Y(Tag2[104]) );
  OAI2B2X1 U1014 ( .A1N(Tag2[103]), .A0(n97), .B0(n1110), .B1(n130), .Y(n7805)
         );
  CLKINVX1 U1015 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[103]), .Y(n1110)
         );
  XOR2X1 U1016 ( .A(n1111), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[103]), 
        .Y(Tag2[103]) );
  OAI2B2X1 U1017 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[102]), .A0(n127), 
        .B0(n526), .B1(n109), .Y(n7804) );
  XOR2X1 U1018 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[102]), .B(n1112), 
        .Y(n526) );
  OAI2B2X1 U1019 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[101]), .A0(n128), 
        .B0(n527), .B1(n109), .Y(n7803) );
  XOR2X1 U1020 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[101]), .B(n1113), 
        .Y(n527) );
  OAI2B2X1 U1021 ( .A1N(Tag2[100]), .A0(n97), .B0(n1114), .B1(n129), .Y(n7802)
         );
  CLKINVX1 U1022 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[100]), .Y(n1114)
         );
  XOR2X1 U1023 ( .A(n1115), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[100]), 
        .Y(Tag2[100]) );
  OAI2B2X1 U1024 ( .A1N(Tag2[99]), .A0(n97), .B0(n1116), .B1(n129), .Y(n7801)
         );
  CLKINVX1 U1025 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[99]), .Y(n1116) );
  XOR2X1 U1026 ( .A(n1117), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[99]), .Y(
        Tag2[99]) );
  OAI2B2X1 U1027 ( .A1N(Tag2[98]), .A0(n97), .B0(n1118), .B1(n129), .Y(n7800)
         );
  CLKINVX1 U1028 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[98]), .Y(n1118) );
  XOR2X1 U1029 ( .A(n1119), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[98]), .Y(
        Tag2[98]) );
  OAI2B2X1 U1030 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[97]), .A0(n128), 
        .B0(n487), .B1(n110), .Y(n7799) );
  XOR2X1 U1031 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[97]), .B(n1120), .Y(
        n487) );
  OAI2B2X1 U1032 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[96]), .A0(n128), 
        .B0(n488), .B1(n109), .Y(n7798) );
  XOR2X1 U1033 ( .A(n1121), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[96]), .Y(
        n488) );
  OAI2B2X1 U1034 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[95]), .A0(n129), 
        .B0(n489), .B1(n110), .Y(n7797) );
  XOR2X1 U1035 ( .A(n1122), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[95]), .Y(
        n489) );
  OAI2B2X1 U1036 ( .A1N(Tag2[94]), .A0(n97), .B0(n1123), .B1(n132), .Y(n7796)
         );
  CLKINVX1 U1037 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[94]), .Y(n1123) );
  XNOR2X1 U1038 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[94]), .B(n1124), 
        .Y(Tag2[94]) );
  OAI2B2X1 U1039 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[93]), .A0(n126), 
        .B0(n490), .B1(n110), .Y(n7795) );
  XOR2X1 U1040 ( .A(n1125), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[93]), .Y(
        n490) );
  OAI2B2X1 U1041 ( .A1N(Tag2[92]), .A0(n97), .B0(n1126), .B1(n132), .Y(n7794)
         );
  CLKINVX1 U1042 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[92]), .Y(n1126) );
  XNOR2X1 U1043 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[92]), .B(n1127), 
        .Y(Tag2[92]) );
  OAI2B2X1 U1044 ( .A1N(Tag2[91]), .A0(n97), .B0(n1128), .B1(n131), .Y(n7793)
         );
  CLKINVX1 U1045 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[91]), .Y(n1128) );
  XOR2X1 U1046 ( .A(n1129), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[91]), .Y(
        Tag2[91]) );
  OAI2B2X1 U1047 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[90]), .A0(n126), 
        .B0(n491), .B1(n110), .Y(n7792) );
  XOR2X1 U1048 ( .A(n1130), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[90]), .Y(
        n491) );
  OAI2B2X1 U1049 ( .A1N(Tag2[89]), .A0(n97), .B0(n1131), .B1(n131), .Y(n7791)
         );
  CLKINVX1 U1050 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[89]), .Y(n1131) );
  XOR2X1 U1051 ( .A(n1132), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[89]), .Y(
        Tag2[89]) );
  OAI2B2X1 U1052 ( .A1N(Tag2[88]), .A0(n97), .B0(n1133), .B1(n130), .Y(n7790)
         );
  CLKINVX1 U1053 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[88]), .Y(n1133) );
  XNOR2X1 U1054 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[88]), .B(n1134), 
        .Y(Tag2[88]) );
  OAI2B2X1 U1055 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[87]), .A0(n126), 
        .B0(n492), .B1(n110), .Y(n7789) );
  XOR2X1 U1056 ( .A(n1135), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[87]), .Y(
        n492) );
  OAI2B2X1 U1057 ( .A1N(Tag2[86]), .A0(n97), .B0(n1136), .B1(n130), .Y(n7788)
         );
  CLKINVX1 U1058 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[86]), .Y(n1136) );
  XNOR2X1 U1059 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[86]), .B(n1137), 
        .Y(Tag2[86]) );
  OAI2B2X1 U1060 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[85]), .A0(n126), 
        .B0(n493), .B1(n110), .Y(n7787) );
  XOR2X1 U1061 ( .A(n1138), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[85]), .Y(
        n493) );
  OAI2B2X1 U1062 ( .A1N(Tag2[84]), .A0(n97), .B0(n1139), .B1(n130), .Y(n7786)
         );
  CLKINVX1 U1063 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[84]), .Y(n1139) );
  XNOR2X1 U1064 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[84]), .B(n1140), 
        .Y(Tag2[84]) );
  OAI2B2X1 U1065 ( .A1N(Tag2[83]), .A0(n98), .B0(n1141), .B1(n130), .Y(n7785)
         );
  CLKINVX1 U1066 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[83]), .Y(n1141) );
  XOR2X1 U1067 ( .A(n1142), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[83]), .Y(
        Tag2[83]) );
  OAI2B2X1 U1068 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[82]), .A0(n126), 
        .B0(n494), .B1(n111), .Y(n7784) );
  XOR2X1 U1069 ( .A(n1143), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[82]), .Y(
        n494) );
  OAI2B2X1 U1070 ( .A1N(Tag2[81]), .A0(n98), .B0(n1144), .B1(n130), .Y(n7783)
         );
  CLKINVX1 U1071 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[81]), .Y(n1144) );
  XOR2X1 U1072 ( .A(n1145), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[81]), .Y(
        Tag2[81]) );
  OAI2B2X1 U1073 ( .A1N(Tag2[80]), .A0(n98), .B0(n1146), .B1(n130), .Y(n7782)
         );
  CLKINVX1 U1074 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[80]), .Y(n1146) );
  XNOR2X1 U1075 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[80]), .B(n1147), 
        .Y(Tag2[80]) );
  OAI2B2X1 U1076 ( .A1N(Tag2[79]), .A0(n98), .B0(n1148), .B1(n129), .Y(n7781)
         );
  CLKINVX1 U1077 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[79]), .Y(n1148) );
  XOR2X1 U1078 ( .A(n1149), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[79]), .Y(
        Tag2[79]) );
  OAI2B2X1 U1079 ( .A1N(Tag2[78]), .A0(n98), .B0(n1150), .B1(n129), .Y(n7780)
         );
  CLKINVX1 U1080 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[78]), .Y(n1150) );
  XNOR2X1 U1081 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[78]), .B(n1151), 
        .Y(Tag2[78]) );
  OAI2B2X1 U1082 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[77]), .A0(n125), 
        .B0(n495), .B1(n111), .Y(n7779) );
  XOR2X1 U1083 ( .A(n1152), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[77]), .Y(
        n495) );
  OAI2B2X1 U1084 ( .A1N(Tag2[76]), .A0(n98), .B0(n1153), .B1(n129), .Y(n7778)
         );
  CLKINVX1 U1085 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[76]), .Y(n1153) );
  XNOR2X1 U1086 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[76]), .B(n1154), 
        .Y(Tag2[76]) );
  OAI2B2X1 U1087 ( .A1N(Tag2[75]), .A0(n98), .B0(n1155), .B1(n129), .Y(n7777)
         );
  CLKINVX1 U1088 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[75]), .Y(n1155) );
  XOR2X1 U1089 ( .A(n1156), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[75]), .Y(
        Tag2[75]) );
  OAI2B2X1 U1090 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[74]), .A0(n125), 
        .B0(n496), .B1(n111), .Y(n7776) );
  XOR2X1 U1091 ( .A(n1157), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[74]), .Y(
        n496) );
  OAI2B2X1 U1092 ( .A1N(Tag2[73]), .A0(n98), .B0(n1158), .B1(n129), .Y(n7775)
         );
  CLKINVX1 U1093 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[73]), .Y(n1158) );
  XOR2X1 U1094 ( .A(n1159), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[73]), .Y(
        Tag2[73]) );
  OAI2B2X1 U1095 ( .A1N(Tag2[72]), .A0(n98), .B0(n1160), .B1(n129), .Y(n7774)
         );
  CLKINVX1 U1096 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[72]), .Y(n1160) );
  XNOR2X1 U1097 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[72]), .B(n1161), 
        .Y(Tag2[72]) );
  OAI2B2X1 U1098 ( .A1N(Tag2[71]), .A0(n98), .B0(n1162), .B1(n129), .Y(n7773)
         );
  CLKINVX1 U1099 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[71]), .Y(n1162) );
  XOR2X1 U1100 ( .A(n1163), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[71]), .Y(
        Tag2[71]) );
  OAI2B2X1 U1101 ( .A1N(Tag2[70]), .A0(n98), .B0(n1164), .B1(n129), .Y(n7772)
         );
  CLKINVX1 U1102 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[70]), .Y(n1164) );
  XNOR2X1 U1103 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[70]), .B(n1165), 
        .Y(Tag2[70]) );
  OAI2B2X1 U1104 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[69]), .A0(n125), 
        .B0(n498), .B1(n111), .Y(n7771) );
  XOR2X1 U1105 ( .A(n1166), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[69]), .Y(
        n498) );
  OAI2B2X1 U1106 ( .A1N(Tag2[68]), .A0(n98), .B0(n1167), .B1(n129), .Y(n7770)
         );
  CLKINVX1 U1107 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[68]), .Y(n1167) );
  XNOR2X1 U1108 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[68]), .B(n1168), 
        .Y(Tag2[68]) );
  OAI2B2X1 U1109 ( .A1N(Tag2[67]), .A0(n98), .B0(n1169), .B1(n130), .Y(n7769)
         );
  CLKINVX1 U1110 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[67]), .Y(n1169) );
  XOR2X1 U1111 ( .A(n1170), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[67]), .Y(
        Tag2[67]) );
  OAI2B2X1 U1112 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[66]), .A0(n125), 
        .B0(n499), .B1(n112), .Y(n7768) );
  XOR2X1 U1113 ( .A(n1171), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[66]), .Y(
        n499) );
  OAI2B2X1 U1114 ( .A1N(Tag2[65]), .A0(n99), .B0(n1172), .B1(n129), .Y(n7767)
         );
  CLKINVX1 U1115 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[65]), .Y(n1172) );
  XOR2X1 U1116 ( .A(n1173), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[65]), .Y(
        Tag2[65]) );
  OAI2B2X1 U1117 ( .A1N(Tag2[64]), .A0(n99), .B0(n1174), .B1(n130), .Y(n7766)
         );
  CLKINVX1 U1118 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[64]), .Y(n1174) );
  XNOR2X1 U1119 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[64]), .B(n1175), 
        .Y(Tag2[64]) );
  OAI2B2X1 U1120 ( .A1N(Tag2[63]), .A0(n99), .B0(n1176), .B1(n129), .Y(n7765)
         );
  CLKINVX1 U1121 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[63]), .Y(n1176) );
  XOR2X1 U1122 ( .A(n1177), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[63]), .Y(
        Tag2[63]) );
  OAI2B2X1 U1123 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[62]), .A0(n124), 
        .B0(n500), .B1(n112), .Y(n7764) );
  XOR2X1 U1124 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[62]), .B(n1178), .Y(
        n500) );
  OAI2B2X1 U1125 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[61]), .A0(n124), 
        .B0(n501), .B1(n112), .Y(n7763) );
  XOR2X1 U1126 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[61]), .B(n1179), .Y(
        n501) );
  OAI2B2X1 U1127 ( .A1N(Tag2[60]), .A0(n99), .B0(n1180), .B1(n130), .Y(n7762)
         );
  CLKINVX1 U1128 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[60]), .Y(n1180) );
  XOR2X1 U1129 ( .A(n1181), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[60]), .Y(
        Tag2[60]) );
  OAI2B2X1 U1130 ( .A1N(Tag2[59]), .A0(n99), .B0(n1182), .B1(n130), .Y(n7761)
         );
  CLKINVX1 U1131 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[59]), .Y(n1182) );
  XOR2X1 U1132 ( .A(n1183), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[59]), .Y(
        Tag2[59]) );
  OAI2B2X1 U1133 ( .A1N(Tag2[58]), .A0(n99), .B0(n1184), .B1(n130), .Y(n7760)
         );
  CLKINVX1 U1134 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[58]), .Y(n1184) );
  XOR2X1 U1135 ( .A(n1185), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[58]), .Y(
        Tag2[58]) );
  OAI2B2X1 U1136 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[57]), .A0(n124), 
        .B0(n502), .B1(n112), .Y(n7759) );
  XOR2X1 U1137 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[57]), .B(n1186), .Y(
        n502) );
  OAI2B2X1 U1138 ( .A1N(Tag2[56]), .A0(n99), .B0(n1187), .B1(n131), .Y(n7758)
         );
  CLKINVX1 U1139 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[56]), .Y(n1187) );
  XOR2X1 U1140 ( .A(n1188), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[56]), .Y(
        Tag2[56]) );
  OAI2B2X1 U1141 ( .A1N(Tag2[55]), .A0(n99), .B0(n1189), .B1(n131), .Y(n7757)
         );
  CLKINVX1 U1142 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[55]), .Y(n1189) );
  XOR2X1 U1143 ( .A(n1190), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[55]), .Y(
        Tag2[55]) );
  OAI2B2X1 U1144 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[54]), .A0(n123), 
        .B0(n503), .B1(n112), .Y(n7756) );
  XOR2X1 U1145 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[54]), .B(n1191), .Y(
        n503) );
  OAI2B2X1 U1146 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[53]), .A0(n123), 
        .B0(n504), .B1(n113), .Y(n7755) );
  XOR2X1 U1147 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[53]), .B(n1192), .Y(
        n504) );
  OAI2B2X1 U1148 ( .A1N(Tag2[52]), .A0(n99), .B0(n1193), .B1(n131), .Y(n7754)
         );
  CLKINVX1 U1149 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[52]), .Y(n1193) );
  XOR2X1 U1150 ( .A(n1194), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[52]), .Y(
        Tag2[52]) );
  OAI2B2X1 U1151 ( .A1N(Tag2[51]), .A0(n99), .B0(n1195), .B1(n131), .Y(n7753)
         );
  CLKINVX1 U1152 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[51]), .Y(n1195) );
  XOR2X1 U1153 ( .A(n1196), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[51]), .Y(
        Tag2[51]) );
  OAI2B2X1 U1154 ( .A1N(Tag2[50]), .A0(n99), .B0(n1197), .B1(n131), .Y(n7752)
         );
  CLKINVX1 U1155 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[50]), .Y(n1197) );
  XOR2X1 U1156 ( .A(n1198), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[50]), .Y(
        Tag2[50]) );
  OAI2B2X1 U1157 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[49]), .A0(n123), 
        .B0(n505), .B1(n113), .Y(n7751) );
  XOR2X1 U1158 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[49]), .B(n1199), .Y(
        n505) );
  OAI2B2X1 U1159 ( .A1N(Tag2[48]), .A0(n99), .B0(n1200), .B1(n131), .Y(n7750)
         );
  CLKINVX1 U1160 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[48]), .Y(n1200) );
  XOR2X1 U1161 ( .A(n1201), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[48]), .Y(
        Tag2[48]) );
  OAI2B2X1 U1162 ( .A1N(Tag2[47]), .A0(n99), .B0(n1202), .B1(n131), .Y(n7749)
         );
  CLKINVX1 U1163 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[47]), .Y(n1202) );
  XOR2X1 U1164 ( .A(n1203), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[47]), .Y(
        Tag2[47]) );
  OAI2B2X1 U1165 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[46]), .A0(n123), 
        .B0(n506), .B1(n113), .Y(n7748) );
  XOR2X1 U1166 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[46]), .B(n1204), .Y(
        n506) );
  OAI2B2X1 U1167 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[45]), .A0(n123), 
        .B0(n507), .B1(n113), .Y(n7747) );
  XOR2X1 U1168 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[45]), .B(n1205), .Y(
        n507) );
  OAI2B2X1 U1169 ( .A1N(Tag2[44]), .A0(n100), .B0(n1206), .B1(n131), .Y(n7746)
         );
  CLKINVX1 U1170 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[44]), .Y(n1206) );
  XOR2X1 U1171 ( .A(n1207), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[44]), .Y(
        Tag2[44]) );
  OAI2B2X1 U1172 ( .A1N(Tag2[43]), .A0(n100), .B0(n1208), .B1(n132), .Y(n7745)
         );
  CLKINVX1 U1173 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[43]), .Y(n1208) );
  XOR2X1 U1174 ( .A(n1209), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[43]), .Y(
        Tag2[43]) );
  OAI2B2X1 U1175 ( .A1N(Tag2[42]), .A0(n100), .B0(n1210), .B1(n131), .Y(n7744)
         );
  CLKINVX1 U1176 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[42]), .Y(n1210) );
  XOR2X1 U1177 ( .A(n1211), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[42]), .Y(
        Tag2[42]) );
  OAI2B2X1 U1178 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[41]), .A0(n123), 
        .B0(n508), .B1(n113), .Y(n7743) );
  XOR2X1 U1179 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[41]), .B(n1212), .Y(
        n508) );
  OAI2B2X1 U1180 ( .A1N(Tag2[40]), .A0(n100), .B0(n1213), .B1(n132), .Y(n7742)
         );
  CLKINVX1 U1181 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[40]), .Y(n1213) );
  XOR2X1 U1182 ( .A(n1214), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[40]), .Y(
        Tag2[40]) );
  OAI2B2X1 U1183 ( .A1N(Tag2[39]), .A0(n100), .B0(n1215), .B1(n132), .Y(n7741)
         );
  CLKINVX1 U1184 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[39]), .Y(n1215) );
  XOR2X1 U1185 ( .A(n1216), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[39]), .Y(
        Tag2[39]) );
  OAI2B2X1 U1186 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[38]), .A0(n123), 
        .B0(n509), .B1(n114), .Y(n7740) );
  XOR2X1 U1187 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[38]), .B(n1217), .Y(
        n509) );
  OAI2B2X1 U1188 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[37]), .A0(n123), 
        .B0(n510), .B1(n114), .Y(n7739) );
  XOR2X1 U1189 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[37]), .B(n1218), .Y(
        n510) );
  OAI2B2X1 U1190 ( .A1N(Tag2[36]), .A0(n100), .B0(n1219), .B1(n132), .Y(n7738)
         );
  CLKINVX1 U1191 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[36]), .Y(n1219) );
  XOR2X1 U1192 ( .A(n1220), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[36]), .Y(
        Tag2[36]) );
  OAI2B2X1 U1193 ( .A1N(Tag2[35]), .A0(n100), .B0(n1221), .B1(n132), .Y(n7737)
         );
  CLKINVX1 U1194 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[35]), .Y(n1221) );
  XOR2X1 U1195 ( .A(n1222), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[35]), .Y(
        Tag2[35]) );
  OAI2B2X1 U1196 ( .A1N(Tag2[34]), .A0(n100), .B0(n1223), .B1(n132), .Y(n7736)
         );
  CLKINVX1 U1197 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[34]), .Y(n1223) );
  XOR2X1 U1198 ( .A(n1224), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[34]), .Y(
        Tag2[34]) );
  OAI2B2X1 U1199 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[33]), .A0(n123), 
        .B0(n511), .B1(n114), .Y(n7735) );
  XOR2X1 U1200 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[33]), .B(n1225), .Y(
        n511) );
  OAI2B2X1 U1201 ( .A1N(Tag2[32]), .A0(n100), .B0(n1226), .B1(n132), .Y(n7734)
         );
  CLKINVX1 U1202 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[32]), .Y(n1226) );
  XOR2X1 U1203 ( .A(n1227), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[32]), .Y(
        Tag2[32]) );
  OAI2B2X1 U1204 ( .A1N(Tag2[31]), .A0(n100), .B0(n1228), .B1(n132), .Y(n7733)
         );
  CLKINVX1 U1205 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[31]), .Y(n1228) );
  XOR2X1 U1206 ( .A(n1229), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[31]), .Y(
        Tag2[31]) );
  OAI2B2X1 U1207 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[30]), .A0(n126), 
        .B0(n512), .B1(n114), .Y(n7732) );
  XOR2X1 U1208 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[30]), .B(n1230), .Y(
        n512) );
  OAI2B2X1 U1209 ( .A1N(Tag2[29]), .A0(n100), .B0(n1231), .B1(n132), .Y(n7731)
         );
  CLKINVX1 U1210 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[29]), .Y(n1231) );
  XOR2X1 U1211 ( .A(n1232), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[29]), .Y(
        Tag2[29]) );
  OAI2B2X1 U1212 ( .A1N(Tag2[28]), .A0(n100), .B0(n1233), .B1(n132), .Y(n7730)
         );
  CLKINVX1 U1213 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[28]), .Y(n1233) );
  XNOR2X1 U1214 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[28]), .B(n1234), 
        .Y(Tag2[28]) );
  OAI2B2X1 U1215 ( .A1N(Tag2[27]), .A0(n100), .B0(n1235), .B1(n132), .Y(n7729)
         );
  CLKINVX1 U1216 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[27]), .Y(n1235) );
  XOR2X1 U1217 ( .A(n1236), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[27]), .Y(
        Tag2[27]) );
  OAI2B2X1 U1218 ( .A1N(Tag2[26]), .A0(n101), .B0(n1237), .B1(n132), .Y(n7728)
         );
  CLKINVX1 U1219 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[26]), .Y(n1237) );
  XOR2X1 U1220 ( .A(n1238), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[26]), .Y(
        Tag2[26]) );
  OAI2B2X1 U1221 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[25]), .A0(n123), 
        .B0(n513), .B1(n114), .Y(n7727) );
  XOR2X1 U1222 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[25]), .B(n1239), .Y(
        n513) );
  OAI2B2X1 U1223 ( .A1N(Tag2[24]), .A0(n101), .B0(n1240), .B1(n132), .Y(n7726)
         );
  CLKINVX1 U1224 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[24]), .Y(n1240) );
  XNOR2X1 U1225 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[24]), .B(n1241), 
        .Y(Tag2[24]) );
  OAI2B2X1 U1226 ( .A1N(Tag2[23]), .A0(n101), .B0(n1242), .B1(n133), .Y(n7725)
         );
  CLKINVX1 U1227 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[23]), .Y(n1242) );
  XOR2X1 U1228 ( .A(n1243), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[23]), .Y(
        Tag2[23]) );
  OAI2B2X1 U1229 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[22]), .A0(n123), 
        .B0(n514), .B1(n114), .Y(n7724) );
  XOR2X1 U1230 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[22]), .B(n1244), .Y(
        n514) );
  OAI2B2X1 U1231 ( .A1N(Tag2[21]), .A0(n101), .B0(n1245), .B1(n133), .Y(n7723)
         );
  CLKINVX1 U1232 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[21]), .Y(n1245) );
  XOR2X1 U1233 ( .A(n1246), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[21]), .Y(
        Tag2[21]) );
  OAI2B2X1 U1234 ( .A1N(Tag2[20]), .A0(n101), .B0(n1247), .B1(n133), .Y(n7722)
         );
  CLKINVX1 U1235 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[20]), .Y(n1247) );
  XNOR2X1 U1236 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[20]), .B(n1248), 
        .Y(Tag2[20]) );
  OAI2B2X1 U1237 ( .A1N(Tag2[19]), .A0(n101), .B0(n1249), .B1(n133), .Y(n7721)
         );
  CLKINVX1 U1238 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[19]), .Y(n1249) );
  XOR2X1 U1239 ( .A(n1250), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[19]), .Y(
        Tag2[19]) );
  OAI2B2X1 U1240 ( .A1N(Tag2[18]), .A0(n101), .B0(n1251), .B1(n133), .Y(n7720)
         );
  CLKINVX1 U1241 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[18]), .Y(n1251) );
  XOR2X1 U1242 ( .A(n1252), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[18]), .Y(
        Tag2[18]) );
  OAI2B2X1 U1243 ( .A1N(Tag2[17]), .A0(n101), .B0(n1253), .B1(n133), .Y(n7719)
         );
  CLKINVX1 U1244 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[17]), .Y(n1253) );
  XOR2X1 U1245 ( .A(n1254), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[17]), .Y(
        Tag2[17]) );
  OAI2B2X1 U1246 ( .A1N(Tag2[16]), .A0(n101), .B0(n1255), .B1(n133), .Y(n7718)
         );
  CLKINVX1 U1247 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[16]), .Y(n1255) );
  XNOR2X1 U1248 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[16]), .B(n1256), 
        .Y(Tag2[16]) );
  OAI2B2X1 U1249 ( .A1N(Tag2[15]), .A0(n101), .B0(n1257), .B1(n133), .Y(n7717)
         );
  CLKINVX1 U1250 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[15]), .Y(n1257) );
  XOR2X1 U1251 ( .A(n1258), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[15]), .Y(
        Tag2[15]) );
  OAI2B2X1 U1252 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[14]), .A0(n123), 
        .B0(n516), .B1(n108), .Y(n7716) );
  XOR2X1 U1253 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[14]), .B(n1259), .Y(
        n516) );
  OAI2B2X1 U1254 ( .A1N(Tag2[13]), .A0(n101), .B0(n1260), .B1(n133), .Y(n7715)
         );
  CLKINVX1 U1255 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[13]), .Y(n1260) );
  XOR2X1 U1256 ( .A(n1261), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[13]), .Y(
        Tag2[13]) );
  OAI2B2X1 U1257 ( .A1N(Tag2[12]), .A0(n101), .B0(n1262), .B1(n133), .Y(n7714)
         );
  CLKINVX1 U1258 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[12]), .Y(n1262) );
  XNOR2X1 U1259 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[12]), .B(n1263), 
        .Y(Tag2[12]) );
  OAI2B2X1 U1260 ( .A1N(Tag2[11]), .A0(n101), .B0(n1264), .B1(n133), .Y(n7713)
         );
  CLKINVX1 U1261 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[11]), .Y(n1264) );
  XOR2X1 U1262 ( .A(n1265), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[11]), .Y(
        Tag2[11]) );
  OAI2B2X1 U1263 ( .A1N(Tag2[10]), .A0(n102), .B0(n1266), .B1(n133), .Y(n7712)
         );
  CLKINVX1 U1264 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[10]), .Y(n1266) );
  XOR2X1 U1265 ( .A(n1267), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[10]), .Y(
        Tag2[10]) );
  OAI2B2X1 U1266 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[9]), .A0(n123), 
        .B0(n486), .B1(n114), .Y(n7711) );
  XOR2X1 U1267 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[9]), .B(n1268), .Y(
        n486) );
  OAI2B2X1 U1268 ( .A1N(Tag2[8]), .A0(n102), .B0(n1269), .B1(n133), .Y(n7710)
         );
  CLKINVX1 U1269 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[8]), .Y(n1269) );
  XNOR2X1 U1270 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[8]), .B(n1270), .Y(
        Tag2[8]) );
  OAI2B2X1 U1271 ( .A1N(Tag2[7]), .A0(n102), .B0(n1271), .B1(n133), .Y(n7709)
         );
  CLKINVX1 U1272 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[7]), .Y(n1271) );
  XOR2X1 U1273 ( .A(n1272), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[7]), .Y(
        Tag2[7]) );
  OAI2B2X1 U1274 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[6]), .A0(n123), 
        .B0(n497), .B1(n114), .Y(n7708) );
  XOR2X1 U1275 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[6]), .B(n1273), .Y(
        n497) );
  OAI2B2X1 U1276 ( .A1N(Tag2[5]), .A0(n102), .B0(n1274), .B1(n133), .Y(n7707)
         );
  CLKINVX1 U1277 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[5]), .Y(n1274) );
  XOR2X1 U1278 ( .A(n1275), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[5]), .Y(
        Tag2[5]) );
  OAI2B2X1 U1279 ( .A1N(Tag2[4]), .A0(n102), .B0(n1276), .B1(n133), .Y(n7706)
         );
  CLKINVX1 U1280 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[4]), .Y(n1276) );
  XNOR2X1 U1281 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[4]), .B(n1277), .Y(
        Tag2[4]) );
  OAI2B2X1 U1282 ( .A1N(Tag2[3]), .A0(n102), .B0(n1278), .B1(n133), .Y(n7705)
         );
  CLKINVX1 U1283 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[3]), .Y(n1278) );
  XOR2X1 U1284 ( .A(n1279), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[3]), .Y(
        Tag2[3]) );
  OAI2B2X1 U1285 ( .A1N(Tag2[2]), .A0(n102), .B0(n1280), .B1(n133), .Y(n7704)
         );
  CLKINVX1 U1286 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[2]), .Y(n1280) );
  XOR2X1 U1287 ( .A(n1281), .B(Inst_forkAE_MainPart2_Auth_Reg_Output[2]), .Y(
        Tag2[2]) );
  OAI2B2X1 U1288 ( .A1N(Inst_forkAE_MainPart2_Auth_Reg_Output[1]), .A0(n123), 
        .B0(n515), .B1(n113), .Y(n7703) );
  XOR2X1 U1289 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[1]), .B(n1282), .Y(
        n515) );
  OAI2B2X1 U1290 ( .A1N(Tag2[0]), .A0(n102), .B0(n1283), .B1(n134), .Y(n7702)
         );
  CLKINVX1 U1291 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[0]), .Y(n1283) );
  XNOR2X1 U1292 ( .A(Inst_forkAE_MainPart2_Auth_Reg_Output[0]), .B(n1284), .Y(
        Tag2[0]) );
  MXI2X1 U1293 ( .A(n1285), .B(n1286), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_127_), .Y(n7445) );
  AOI21X1 U1294 ( .A0(n1287), .A1(n41), .B0(n66), .Y(n1286) );
  CLKNAND2X2 U1295 ( .A(n23), .B(n1288), .Y(n1285) );
  MXI2X1 U1296 ( .A(n1289), .B(n1290), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_126_), .Y(n7444) );
  AOI21X1 U1297 ( .A0(n1291), .A1(n41), .B0(n65), .Y(n1290) );
  NAND2BX1 U1298 ( .AN(n1291), .B(n34), .Y(n1289) );
  MXI2X1 U1299 ( .A(n1292), .B(n1293), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_125_), .Y(n7443) );
  AOI21X1 U1300 ( .A0(n1294), .A1(n41), .B0(n65), .Y(n1293) );
  NAND2BX1 U1301 ( .AN(n1294), .B(n33), .Y(n1292) );
  MXI2X1 U1302 ( .A(n1295), .B(n1296), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_124_), .Y(n7442) );
  AOI21X1 U1303 ( .A0(n1297), .A1(n41), .B0(n65), .Y(n1296) );
  NAND2BX1 U1304 ( .AN(n1297), .B(n33), .Y(n1295) );
  MXI2X1 U1305 ( .A(n1298), .B(n1299), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_123_), .Y(n7441) );
  AOI21X1 U1306 ( .A0(n1300), .A1(n41), .B0(n65), .Y(n1299) );
  NAND2BX1 U1307 ( .AN(n1300), .B(n33), .Y(n1298) );
  MXI2X1 U1308 ( .A(n1301), .B(n1302), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_122_), .Y(n7440) );
  AOI21X1 U1309 ( .A0(n1303), .A1(n44), .B0(n65), .Y(n1302) );
  NAND2BX1 U1310 ( .AN(n1303), .B(n34), .Y(n1301) );
  MXI2X1 U1311 ( .A(n1304), .B(n1305), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_121_), .Y(n7439) );
  AOI21X1 U1312 ( .A0(n1306), .A1(n35), .B0(n65), .Y(n1305) );
  NAND2BX1 U1313 ( .AN(n1306), .B(n33), .Y(n1304) );
  MXI2X1 U1314 ( .A(n1307), .B(n1308), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_120_), .Y(n7438) );
  AOI21X1 U1315 ( .A0(n1309), .A1(n41), .B0(n65), .Y(n1308) );
  NAND2BX1 U1316 ( .AN(n1309), .B(n34), .Y(n1307) );
  MXI2X1 U1317 ( .A(n1310), .B(n1311), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_119_), .Y(n7437) );
  AOI2B1X1 U1318 ( .A1N(n1312), .A0(n32), .B0(n83), .Y(n1311) );
  CLKNAND2X2 U1319 ( .A(n22), .B(n1312), .Y(n1310) );
  MXI2X1 U1320 ( .A(n1313), .B(n1314), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_118_), .Y(n7436) );
  AOI21X1 U1321 ( .A0(n1315), .A1(n42), .B0(n65), .Y(n1314) );
  CLKNAND2X2 U1322 ( .A(n22), .B(n1316), .Y(n1313) );
  MXI2X1 U1323 ( .A(n1317), .B(n1318), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_117_), .Y(n7435) );
  AOI21X1 U1324 ( .A0(n1319), .A1(n42), .B0(n65), .Y(n1318) );
  CLKNAND2X2 U1325 ( .A(n22), .B(n1320), .Y(n1317) );
  MXI2X1 U1326 ( .A(n1321), .B(n1322), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_116_), .Y(n7434) );
  AOI21X1 U1327 ( .A0(n1323), .A1(n42), .B0(n65), .Y(n1322) );
  CLKNAND2X2 U1328 ( .A(n22), .B(n1324), .Y(n1321) );
  MXI2X1 U1329 ( .A(n1325), .B(n1326), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_115_), .Y(n7433) );
  AOI21X1 U1330 ( .A0(n1327), .A1(n42), .B0(n65), .Y(n1326) );
  CLKNAND2X2 U1331 ( .A(n22), .B(n1328), .Y(n1325) );
  MXI2X1 U1332 ( .A(n1329), .B(n1330), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_114_), .Y(n7432) );
  AOI21X1 U1333 ( .A0(n1331), .A1(n42), .B0(n69), .Y(n1330) );
  CLKNAND2X2 U1334 ( .A(n22), .B(n1332), .Y(n1329) );
  MXI2X1 U1335 ( .A(n1333), .B(n1334), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_113_), .Y(n7431) );
  AOI21X1 U1336 ( .A0(n1335), .A1(n42), .B0(n82), .Y(n1334) );
  CLKNAND2X2 U1337 ( .A(n21), .B(n1336), .Y(n1333) );
  MXI2X1 U1338 ( .A(n1337), .B(n1338), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_112_), .Y(n7430) );
  AOI21X1 U1339 ( .A0(n1339), .A1(n42), .B0(n82), .Y(n1338) );
  CLKNAND2X2 U1340 ( .A(n21), .B(n1340), .Y(n1337) );
  MXI2X1 U1341 ( .A(n1341), .B(n1342), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_111_), .Y(n7429) );
  AOI2B1X1 U1342 ( .A1N(n1343), .A0(n32), .B0(n83), .Y(n1342) );
  CLKNAND2X2 U1343 ( .A(n21), .B(n1343), .Y(n1341) );
  MXI2X1 U1344 ( .A(n1344), .B(n1345), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_110_), .Y(n7428) );
  AOI21X1 U1345 ( .A0(n1346), .A1(n42), .B0(n82), .Y(n1345) );
  CLKNAND2X2 U1346 ( .A(n21), .B(n1347), .Y(n1344) );
  MXI2X1 U1347 ( .A(n1348), .B(n1349), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_109_), .Y(n7427) );
  AOI21X1 U1348 ( .A0(n1350), .A1(n42), .B0(n82), .Y(n1349) );
  CLKNAND2X2 U1349 ( .A(n21), .B(n1351), .Y(n1348) );
  MXI2X1 U1350 ( .A(n1352), .B(n1353), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_108_), .Y(n7426) );
  AOI21X1 U1351 ( .A0(n1354), .A1(n43), .B0(n81), .Y(n1353) );
  CLKNAND2X2 U1352 ( .A(n21), .B(n1355), .Y(n1352) );
  MXI2X1 U1353 ( .A(n1356), .B(n1357), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_107_), .Y(n7425) );
  AOI21X1 U1354 ( .A0(n1358), .A1(n43), .B0(n82), .Y(n1357) );
  CLKNAND2X2 U1355 ( .A(n21), .B(n1359), .Y(n1356) );
  MXI2X1 U1356 ( .A(n1360), .B(n1361), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_106_), .Y(n7424) );
  AOI21X1 U1357 ( .A0(n1362), .A1(n43), .B0(n81), .Y(n1361) );
  CLKNAND2X2 U1358 ( .A(n20), .B(n1363), .Y(n1360) );
  MXI2X1 U1359 ( .A(n1364), .B(n1365), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_105_), .Y(n7423) );
  AOI21X1 U1360 ( .A0(n1366), .A1(n43), .B0(n81), .Y(n1365) );
  CLKNAND2X2 U1361 ( .A(n20), .B(n1367), .Y(n1364) );
  MXI2X1 U1362 ( .A(n1368), .B(n1369), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_104_), .Y(n7422) );
  AOI21X1 U1363 ( .A0(n1370), .A1(n43), .B0(n81), .Y(n1369) );
  CLKNAND2X2 U1364 ( .A(n20), .B(n1371), .Y(n1368) );
  MXI2X1 U1365 ( .A(n1372), .B(n1373), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_103_), .Y(n7421) );
  AOI2B1X1 U1366 ( .A1N(n1374), .A0(n32), .B0(n83), .Y(n1373) );
  CLKNAND2X2 U1367 ( .A(n20), .B(n1374), .Y(n1372) );
  MXI2X1 U1368 ( .A(n1375), .B(n1376), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_102_), .Y(n7420) );
  AOI21X1 U1369 ( .A0(n1377), .A1(n43), .B0(n81), .Y(n1376) );
  CLKNAND2X2 U1370 ( .A(n20), .B(n1378), .Y(n1375) );
  MXI2X1 U1371 ( .A(n1379), .B(n1380), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_101_), .Y(n7419) );
  AOI21X1 U1372 ( .A0(n1381), .A1(n43), .B0(n81), .Y(n1380) );
  CLKNAND2X2 U1373 ( .A(n20), .B(n1382), .Y(n1379) );
  MXI2X1 U1374 ( .A(n1383), .B(n1384), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_100_), .Y(n7418) );
  AOI21X1 U1375 ( .A0(n1385), .A1(n43), .B0(n81), .Y(n1384) );
  CLKNAND2X2 U1376 ( .A(n20), .B(n1386), .Y(n1383) );
  MXI2X1 U1377 ( .A(n1387), .B(n1388), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_99_), .Y(n7417) );
  AOI21X1 U1378 ( .A0(n1389), .A1(n41), .B0(n81), .Y(n1388) );
  CLKNAND2X2 U1379 ( .A(n19), .B(n1390), .Y(n1387) );
  MXI2X1 U1380 ( .A(n1391), .B(n1392), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_98_), .Y(n7416) );
  AOI21X1 U1381 ( .A0(n1393), .A1(n44), .B0(n81), .Y(n1392) );
  CLKNAND2X2 U1382 ( .A(n19), .B(n1394), .Y(n1391) );
  MXI2X1 U1383 ( .A(n1395), .B(n1396), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_97_), .Y(n7415) );
  AOI21X1 U1384 ( .A0(n1397), .A1(n44), .B0(n81), .Y(n1396) );
  CLKNAND2X2 U1385 ( .A(n19), .B(n1398), .Y(n1395) );
  MXI2X1 U1386 ( .A(n1399), .B(n1400), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_96_), .Y(n7414) );
  AOI21X1 U1387 ( .A0(n1401), .A1(n44), .B0(n81), .Y(n1400) );
  CLKNAND2X2 U1388 ( .A(n19), .B(n1402), .Y(n1399) );
  MXI2X1 U1389 ( .A(n1403), .B(n1404), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_95_), .Y(n7413) );
  AOI2B1X1 U1390 ( .A1N(n1405), .A0(n32), .B0(n84), .Y(n1404) );
  CLKNAND2X2 U1391 ( .A(n19), .B(n1405), .Y(n1403) );
  MXI2X1 U1392 ( .A(n1406), .B(n1407), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_94_), .Y(n7412) );
  AOI21X1 U1393 ( .A0(n1408), .A1(n44), .B0(n81), .Y(n1407) );
  CLKNAND2X2 U1394 ( .A(n19), .B(n1409), .Y(n1406) );
  MXI2X1 U1395 ( .A(n1410), .B(n1411), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_93_), .Y(n7411) );
  AOI21X1 U1396 ( .A0(n1412), .A1(n44), .B0(n80), .Y(n1411) );
  CLKNAND2X2 U1397 ( .A(n19), .B(n1413), .Y(n1410) );
  MXI2X1 U1398 ( .A(n1414), .B(n1415), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_92_), .Y(n7410) );
  AOI21X1 U1399 ( .A0(n1416), .A1(n44), .B0(n80), .Y(n1415) );
  CLKNAND2X2 U1400 ( .A(n18), .B(n1417), .Y(n1414) );
  MXI2X1 U1401 ( .A(n1418), .B(n1419), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_91_), .Y(n7409) );
  AOI21X1 U1402 ( .A0(n1420), .A1(n44), .B0(n80), .Y(n1419) );
  CLKNAND2X2 U1403 ( .A(n18), .B(n1421), .Y(n1418) );
  MXI2X1 U1404 ( .A(n1422), .B(n1423), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_90_), .Y(n7408) );
  AOI21X1 U1405 ( .A0(n1424), .A1(n44), .B0(n80), .Y(n1423) );
  CLKNAND2X2 U1406 ( .A(n18), .B(n1425), .Y(n1422) );
  MXI2X1 U1407 ( .A(n1426), .B(n1427), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_89_), .Y(n7407) );
  AOI21X1 U1408 ( .A0(n1428), .A1(n44), .B0(n80), .Y(n1427) );
  CLKNAND2X2 U1409 ( .A(n18), .B(n1429), .Y(n1426) );
  MXI2X1 U1410 ( .A(n1430), .B(n1431), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_88_), .Y(n7406) );
  AOI21X1 U1411 ( .A0(n1432), .A1(n45), .B0(n80), .Y(n1431) );
  CLKNAND2X2 U1412 ( .A(n18), .B(n1433), .Y(n1430) );
  MXI2X1 U1413 ( .A(n1434), .B(n1435), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_87_), .Y(n7405) );
  AOI2B1X1 U1414 ( .A1N(n1436), .A0(n33), .B0(n84), .Y(n1435) );
  CLKNAND2X2 U1415 ( .A(n18), .B(n1436), .Y(n1434) );
  MXI2X1 U1416 ( .A(n1437), .B(n1438), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_86_), .Y(n7404) );
  AOI21X1 U1417 ( .A0(n1439), .A1(n45), .B0(n80), .Y(n1438) );
  CLKNAND2X2 U1418 ( .A(n17), .B(n1440), .Y(n1437) );
  MXI2X1 U1419 ( .A(n1441), .B(n1442), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_85_), .Y(n7403) );
  AOI21X1 U1420 ( .A0(n1443), .A1(n45), .B0(n80), .Y(n1442) );
  CLKNAND2X2 U1421 ( .A(n17), .B(n1444), .Y(n1441) );
  MXI2X1 U1422 ( .A(n1445), .B(n1446), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_84_), .Y(n7402) );
  AOI21X1 U1423 ( .A0(n1447), .A1(n45), .B0(n80), .Y(n1446) );
  CLKNAND2X2 U1424 ( .A(n17), .B(n1448), .Y(n1445) );
  MXI2X1 U1425 ( .A(n1449), .B(n1450), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_83_), .Y(n7401) );
  AOI21X1 U1426 ( .A0(n1451), .A1(n45), .B0(n80), .Y(n1450) );
  CLKNAND2X2 U1427 ( .A(n17), .B(n1452), .Y(n1449) );
  MXI2X1 U1428 ( .A(n1453), .B(n1454), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_82_), .Y(n7400) );
  AOI21X1 U1429 ( .A0(n1455), .A1(n45), .B0(n80), .Y(n1454) );
  CLKNAND2X2 U1430 ( .A(n17), .B(n1456), .Y(n1453) );
  MXI2X1 U1431 ( .A(n1457), .B(n1458), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_81_), .Y(n7399) );
  AOI21X1 U1432 ( .A0(n1459), .A1(n45), .B0(n79), .Y(n1458) );
  CLKNAND2X2 U1433 ( .A(n17), .B(n1460), .Y(n1457) );
  MXI2X1 U1434 ( .A(n1461), .B(n1462), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_80_), .Y(n7398) );
  AOI21X1 U1435 ( .A0(n1463), .A1(n45), .B0(n79), .Y(n1462) );
  CLKNAND2X2 U1436 ( .A(n17), .B(n1464), .Y(n1461) );
  MXI2X1 U1437 ( .A(n1465), .B(n1466), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_79_), .Y(n7397) );
  AOI2B1X1 U1438 ( .A1N(n1467), .A0(n32), .B0(n84), .Y(n1466) );
  CLKNAND2X2 U1439 ( .A(n16), .B(n1467), .Y(n1465) );
  MXI2X1 U1440 ( .A(n1468), .B(n1469), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_78_), .Y(n7396) );
  AOI21X1 U1441 ( .A0(n1470), .A1(n46), .B0(n79), .Y(n1469) );
  CLKNAND2X2 U1442 ( .A(n16), .B(n1471), .Y(n1468) );
  MXI2X1 U1443 ( .A(n1472), .B(n1473), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_77_), .Y(n7395) );
  AOI21X1 U1444 ( .A0(n1474), .A1(n46), .B0(n79), .Y(n1473) );
  CLKNAND2X2 U1445 ( .A(n16), .B(n1475), .Y(n1472) );
  MXI2X1 U1446 ( .A(n1476), .B(n1477), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_76_), .Y(n7394) );
  AOI21X1 U1447 ( .A0(n1478), .A1(n46), .B0(n79), .Y(n1477) );
  CLKNAND2X2 U1448 ( .A(n16), .B(n1479), .Y(n1476) );
  MXI2X1 U1449 ( .A(n1480), .B(n1481), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_75_), .Y(n7393) );
  AOI21X1 U1450 ( .A0(n1482), .A1(n46), .B0(n79), .Y(n1481) );
  CLKNAND2X2 U1451 ( .A(n16), .B(n1483), .Y(n1480) );
  MXI2X1 U1452 ( .A(n1484), .B(n1485), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_74_), .Y(n7392) );
  AOI21X1 U1453 ( .A0(n1486), .A1(n46), .B0(n79), .Y(n1485) );
  CLKNAND2X2 U1454 ( .A(n16), .B(n1487), .Y(n1484) );
  MXI2X1 U1455 ( .A(n1488), .B(n1489), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_73_), .Y(n7391) );
  AOI21X1 U1456 ( .A0(n1490), .A1(n46), .B0(n79), .Y(n1489) );
  CLKNAND2X2 U1457 ( .A(n16), .B(n1491), .Y(n1488) );
  MXI2X1 U1458 ( .A(n1492), .B(n1493), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_72_), .Y(n7390) );
  AOI21X1 U1459 ( .A0(n1494), .A1(n46), .B0(n79), .Y(n1493) );
  CLKNAND2X2 U1460 ( .A(n15), .B(n1495), .Y(n1492) );
  MXI2X1 U1461 ( .A(n1496), .B(n1497), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_71_), .Y(n7389) );
  AOI2B1X1 U1462 ( .A1N(n1498), .A0(n33), .B0(n84), .Y(n1497) );
  CLKNAND2X2 U1463 ( .A(n15), .B(n1498), .Y(n1496) );
  MXI2X1 U1464 ( .A(n1499), .B(n1500), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_70_), .Y(n7388) );
  AOI21X1 U1465 ( .A0(n1501), .A1(n46), .B0(n79), .Y(n1500) );
  CLKNAND2X2 U1466 ( .A(n15), .B(n1502), .Y(n1499) );
  MXI2X1 U1467 ( .A(n1503), .B(n1504), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_69_), .Y(n7387) );
  AOI21X1 U1468 ( .A0(n1505), .A1(n46), .B0(n79), .Y(n1504) );
  CLKNAND2X2 U1469 ( .A(n15), .B(n1506), .Y(n1503) );
  MXI2X1 U1470 ( .A(n1507), .B(n1508), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_68_), .Y(n7386) );
  AOI21X1 U1471 ( .A0(n1509), .A1(n47), .B0(n79), .Y(n1508) );
  CLKNAND2X2 U1472 ( .A(n15), .B(n1510), .Y(n1507) );
  MXI2X1 U1473 ( .A(n1511), .B(n1512), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_67_), .Y(n7385) );
  AOI21X1 U1474 ( .A0(n1513), .A1(n47), .B0(n78), .Y(n1512) );
  CLKNAND2X2 U1475 ( .A(n15), .B(n1514), .Y(n1511) );
  MXI2X1 U1476 ( .A(n1515), .B(n1516), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_66_), .Y(n7384) );
  AOI21X1 U1477 ( .A0(n1517), .A1(n47), .B0(n78), .Y(n1516) );
  CLKNAND2X2 U1478 ( .A(n15), .B(n1518), .Y(n1515) );
  MXI2X1 U1479 ( .A(n1519), .B(n1520), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_65_), .Y(n7383) );
  AOI21X1 U1480 ( .A0(n1521), .A1(n47), .B0(n78), .Y(n1520) );
  CLKNAND2X2 U1481 ( .A(n14), .B(n1522), .Y(n1519) );
  MXI2X1 U1482 ( .A(n1523), .B(n1524), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_64_), .Y(n7382) );
  AOI21X1 U1483 ( .A0(n1525), .A1(n47), .B0(n78), .Y(n1524) );
  CLKNAND2X2 U1484 ( .A(n14), .B(n1526), .Y(n1523) );
  MXI2X1 U1485 ( .A(n1527), .B(n1528), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_63_), .Y(n7381) );
  AOI2B1X1 U1486 ( .A1N(n1529), .A0(n32), .B0(n84), .Y(n1528) );
  CLKNAND2X2 U1487 ( .A(n14), .B(n1529), .Y(n1527) );
  MXI2X1 U1488 ( .A(n1530), .B(n1531), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_62_), .Y(n7380) );
  AOI21X1 U1489 ( .A0(n1532), .A1(n47), .B0(n78), .Y(n1531) );
  CLKNAND2X2 U1490 ( .A(n14), .B(n1533), .Y(n1530) );
  MXI2X1 U1491 ( .A(n1534), .B(n1535), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_61_), .Y(n7379) );
  AOI21X1 U1492 ( .A0(n1536), .A1(n47), .B0(n78), .Y(n1535) );
  CLKNAND2X2 U1493 ( .A(n14), .B(n1537), .Y(n1534) );
  MXI2X1 U1494 ( .A(n1538), .B(n1539), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_60_), .Y(n7378) );
  AOI21X1 U1495 ( .A0(n1540), .A1(n47), .B0(n78), .Y(n1539) );
  CLKNAND2X2 U1496 ( .A(n14), .B(n1541), .Y(n1538) );
  MXI2X1 U1497 ( .A(n1542), .B(n1543), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_59_), .Y(n7377) );
  AOI21X1 U1498 ( .A0(n1544), .A1(n47), .B0(n78), .Y(n1543) );
  CLKNAND2X2 U1499 ( .A(n18), .B(n1545), .Y(n1542) );
  MXI2X1 U1500 ( .A(n1546), .B(n1547), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_58_), .Y(n7376) );
  AOI21X1 U1501 ( .A0(n1548), .A1(n48), .B0(n78), .Y(n1547) );
  CLKNAND2X2 U1502 ( .A(n31), .B(n1549), .Y(n1546) );
  MXI2X1 U1503 ( .A(n1550), .B(n1551), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_57_), .Y(n7375) );
  AOI21X1 U1504 ( .A0(n1552), .A1(n48), .B0(n78), .Y(n1551) );
  CLKNAND2X2 U1505 ( .A(n31), .B(n1553), .Y(n1550) );
  MXI2X1 U1506 ( .A(n1554), .B(n1555), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_56_), .Y(n7374) );
  AOI21X1 U1507 ( .A0(n1556), .A1(n48), .B0(n78), .Y(n1555) );
  CLKNAND2X2 U1508 ( .A(n30), .B(n1557), .Y(n1554) );
  MXI2X1 U1509 ( .A(n1558), .B(n1559), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_55_), .Y(n7373) );
  AOI2B1X1 U1510 ( .A1N(n1560), .A0(n33), .B0(n84), .Y(n1559) );
  CLKNAND2X2 U1511 ( .A(n30), .B(n1560), .Y(n1558) );
  MXI2X1 U1512 ( .A(n1561), .B(n1562), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_54_), .Y(n7372) );
  AOI21X1 U1513 ( .A0(n1563), .A1(n35), .B0(n77), .Y(n1562) );
  CLKNAND2X2 U1514 ( .A(n31), .B(n1564), .Y(n1561) );
  MXI2X1 U1515 ( .A(n1565), .B(n1566), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_53_), .Y(n7371) );
  AOI21X1 U1516 ( .A0(n1567), .A1(n35), .B0(n77), .Y(n1566) );
  CLKNAND2X2 U1517 ( .A(n29), .B(n1568), .Y(n1565) );
  MXI2X1 U1518 ( .A(n1569), .B(n1570), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_52_), .Y(n7370) );
  AOI21X1 U1519 ( .A0(n1571), .A1(n35), .B0(n77), .Y(n1570) );
  CLKNAND2X2 U1520 ( .A(n30), .B(n1572), .Y(n1569) );
  MXI2X1 U1521 ( .A(n1573), .B(n1574), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_51_), .Y(n7369) );
  AOI21X1 U1522 ( .A0(n1575), .A1(n35), .B0(n77), .Y(n1574) );
  CLKNAND2X2 U1523 ( .A(n30), .B(n1576), .Y(n1573) );
  MXI2X1 U1524 ( .A(n1577), .B(n1578), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_50_), .Y(n7368) );
  AOI21X1 U1525 ( .A0(n1579), .A1(n36), .B0(n77), .Y(n1578) );
  CLKNAND2X2 U1526 ( .A(n30), .B(n1580), .Y(n1577) );
  MXI2X1 U1527 ( .A(n1581), .B(n1582), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_49_), .Y(n7367) );
  AOI21X1 U1528 ( .A0(n1583), .A1(n37), .B0(n77), .Y(n1582) );
  CLKNAND2X2 U1529 ( .A(n30), .B(n1584), .Y(n1581) );
  MXI2X1 U1530 ( .A(n1585), .B(n1586), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_48_), .Y(n7366) );
  AOI21X1 U1531 ( .A0(n1587), .A1(n36), .B0(n77), .Y(n1586) );
  CLKNAND2X2 U1532 ( .A(n29), .B(n1588), .Y(n1585) );
  MXI2X1 U1533 ( .A(n1589), .B(n1590), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_47_), .Y(n7365) );
  AOI2B1X1 U1534 ( .A1N(n1591), .A0(n32), .B0(n84), .Y(n1590) );
  CLKNAND2X2 U1535 ( .A(n29), .B(n1591), .Y(n1589) );
  MXI2X1 U1536 ( .A(n1592), .B(n1593), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_46_), .Y(n7364) );
  AOI21X1 U1537 ( .A0(n1594), .A1(n35), .B0(n77), .Y(n1593) );
  CLKNAND2X2 U1538 ( .A(n30), .B(n1595), .Y(n1592) );
  MXI2X1 U1539 ( .A(n1596), .B(n1597), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_45_), .Y(n7363) );
  AOI21X1 U1540 ( .A0(n1598), .A1(n35), .B0(n77), .Y(n1597) );
  CLKNAND2X2 U1541 ( .A(n29), .B(n1599), .Y(n1596) );
  MXI2X1 U1542 ( .A(n1600), .B(n1601), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_44_), .Y(n7362) );
  AOI21X1 U1543 ( .A0(n1602), .A1(n35), .B0(n77), .Y(n1601) );
  CLKNAND2X2 U1544 ( .A(n29), .B(n1603), .Y(n1600) );
  MXI2X1 U1545 ( .A(n1604), .B(n1605), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_43_), .Y(n7361) );
  AOI21X1 U1546 ( .A0(n1606), .A1(n36), .B0(n77), .Y(n1605) );
  CLKNAND2X2 U1547 ( .A(n29), .B(n1607), .Y(n1604) );
  MXI2X1 U1548 ( .A(n1608), .B(n1609), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_42_), .Y(n7360) );
  AOI21X1 U1549 ( .A0(n1610), .A1(n36), .B0(n76), .Y(n1609) );
  CLKNAND2X2 U1550 ( .A(n29), .B(n1611), .Y(n1608) );
  MXI2X1 U1551 ( .A(n1612), .B(n1613), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_41_), .Y(n7359) );
  AOI21X1 U1552 ( .A0(n1614), .A1(n36), .B0(n76), .Y(n1613) );
  CLKNAND2X2 U1553 ( .A(n29), .B(n1615), .Y(n1612) );
  MXI2X1 U1554 ( .A(n1616), .B(n1617), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_40_), .Y(n7358) );
  AOI21X1 U1555 ( .A0(n1618), .A1(n36), .B0(n76), .Y(n1617) );
  CLKNAND2X2 U1556 ( .A(n28), .B(n1619), .Y(n1616) );
  MXI2X1 U1557 ( .A(n1620), .B(n1621), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_39_), .Y(n7357) );
  AOI2B1X1 U1558 ( .A1N(n1622), .A0(n32), .B0(n84), .Y(n1621) );
  CLKNAND2X2 U1559 ( .A(n28), .B(n1622), .Y(n1620) );
  MXI2X1 U1560 ( .A(n1623), .B(n1624), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_38_), .Y(n7356) );
  AOI21X1 U1561 ( .A0(n1625), .A1(n36), .B0(n76), .Y(n1624) );
  CLKNAND2X2 U1562 ( .A(n28), .B(n1626), .Y(n1623) );
  MXI2X1 U1563 ( .A(n1627), .B(n1628), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_37_), .Y(n7355) );
  AOI21X1 U1564 ( .A0(n1629), .A1(n36), .B0(n76), .Y(n1628) );
  CLKNAND2X2 U1565 ( .A(n28), .B(n1630), .Y(n1627) );
  MXI2X1 U1566 ( .A(n1631), .B(n1632), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_36_), .Y(n7354) );
  AOI21X1 U1567 ( .A0(n1633), .A1(n36), .B0(n76), .Y(n1632) );
  CLKNAND2X2 U1568 ( .A(n28), .B(n1634), .Y(n1631) );
  MXI2X1 U1569 ( .A(n1635), .B(n1636), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_35_), .Y(n7353) );
  AOI21X1 U1570 ( .A0(n1637), .A1(n36), .B0(n76), .Y(n1636) );
  CLKNAND2X2 U1571 ( .A(n27), .B(n1638), .Y(n1635) );
  MXI2X1 U1572 ( .A(n1639), .B(n1640), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_34_), .Y(n7352) );
  AOI21X1 U1573 ( .A0(n1641), .A1(n37), .B0(n76), .Y(n1640) );
  CLKNAND2X2 U1574 ( .A(n27), .B(n1642), .Y(n1639) );
  MXI2X1 U1575 ( .A(n1643), .B(n1644), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_33_), .Y(n7351) );
  AOI21X1 U1576 ( .A0(n1645), .A1(n37), .B0(n76), .Y(n1644) );
  CLKNAND2X2 U1577 ( .A(n27), .B(n1646), .Y(n1643) );
  MXI2X1 U1578 ( .A(n1647), .B(n1648), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_32_), .Y(n7350) );
  AOI21X1 U1579 ( .A0(n1649), .A1(n37), .B0(n76), .Y(n1648) );
  CLKNAND2X2 U1580 ( .A(n27), .B(n1650), .Y(n1647) );
  MXI2X1 U1581 ( .A(n1651), .B(n1652), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_31_), .Y(n7349) );
  AOI2B1X1 U1582 ( .A1N(n1653), .A0(n33), .B0(n84), .Y(n1652) );
  CLKNAND2X2 U1583 ( .A(n27), .B(n1653), .Y(n1651) );
  MXI2X1 U1584 ( .A(n1654), .B(n1655), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_30_), .Y(n7348) );
  AOI21X1 U1585 ( .A0(n1656), .A1(n37), .B0(n76), .Y(n1655) );
  CLKNAND2X2 U1586 ( .A(n27), .B(n1657), .Y(n1654) );
  MXI2X1 U1587 ( .A(n1658), .B(n1659), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_29_), .Y(n7347) );
  AOI21X1 U1588 ( .A0(n1660), .A1(n37), .B0(n75), .Y(n1659) );
  CLKNAND2X2 U1589 ( .A(n27), .B(n1661), .Y(n1658) );
  MXI2X1 U1590 ( .A(n1662), .B(n1663), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_28_), .Y(n7346) );
  AOI21X1 U1591 ( .A0(n1664), .A1(n37), .B0(n75), .Y(n1663) );
  CLKNAND2X2 U1592 ( .A(n26), .B(n1665), .Y(n1662) );
  MXI2X1 U1593 ( .A(n1666), .B(n1667), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_27_), .Y(n7345) );
  AOI21X1 U1594 ( .A0(n1668), .A1(n37), .B0(n75), .Y(n1667) );
  CLKNAND2X2 U1595 ( .A(n26), .B(n1669), .Y(n1666) );
  MXI2X1 U1596 ( .A(n1670), .B(n1671), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_26_), .Y(n7344) );
  AOI21X1 U1597 ( .A0(n1672), .A1(n37), .B0(n78), .Y(n1671) );
  CLKNAND2X2 U1598 ( .A(n26), .B(n1673), .Y(n1670) );
  MXI2X1 U1599 ( .A(n1674), .B(n1675), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_25_), .Y(n7343) );
  AOI21X1 U1600 ( .A0(n1676), .A1(n38), .B0(n75), .Y(n1675) );
  CLKNAND2X2 U1601 ( .A(n26), .B(n1677), .Y(n1674) );
  MXI2X1 U1602 ( .A(n1678), .B(n1679), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_24_), .Y(n7342) );
  AOI21X1 U1603 ( .A0(n1680), .A1(n38), .B0(n75), .Y(n1679) );
  CLKNAND2X2 U1604 ( .A(n26), .B(n1681), .Y(n1678) );
  MXI2X1 U1605 ( .A(n1682), .B(n1683), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_23_), .Y(n7341) );
  AOI2B1X1 U1606 ( .A1N(n1684), .A0(n33), .B0(n84), .Y(n1683) );
  CLKNAND2X2 U1607 ( .A(n26), .B(n1684), .Y(n1682) );
  MXI2X1 U1608 ( .A(n1685), .B(n1686), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_22_), .Y(n7340) );
  AOI21X1 U1609 ( .A0(n1687), .A1(n38), .B0(n75), .Y(n1686) );
  CLKNAND2X2 U1610 ( .A(n26), .B(n1688), .Y(n1685) );
  MXI2X1 U1611 ( .A(n1689), .B(n1690), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_21_), .Y(n7339) );
  AOI21X1 U1612 ( .A0(n1691), .A1(n38), .B0(n75), .Y(n1690) );
  CLKNAND2X2 U1613 ( .A(n25), .B(n1692), .Y(n1689) );
  MXI2X1 U1614 ( .A(n1693), .B(n1694), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_20_), .Y(n7338) );
  AOI21X1 U1615 ( .A0(n1695), .A1(n38), .B0(n75), .Y(n1694) );
  CLKNAND2X2 U1616 ( .A(n25), .B(n1696), .Y(n1693) );
  MXI2X1 U1617 ( .A(n1697), .B(n1698), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_19_), .Y(n7337) );
  AOI21X1 U1618 ( .A0(n1699), .A1(n38), .B0(n75), .Y(n1698) );
  CLKNAND2X2 U1619 ( .A(n25), .B(n1700), .Y(n1697) );
  MXI2X1 U1620 ( .A(n1701), .B(n1702), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_18_), .Y(n7336) );
  AOI21X1 U1621 ( .A0(n1703), .A1(n38), .B0(n75), .Y(n1702) );
  CLKNAND2X2 U1622 ( .A(n25), .B(n1704), .Y(n1701) );
  MXI2X1 U1623 ( .A(n1705), .B(n1706), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_17_), .Y(n7335) );
  AOI21X1 U1624 ( .A0(n1707), .A1(n38), .B0(n75), .Y(n1706) );
  CLKNAND2X2 U1625 ( .A(n25), .B(n1708), .Y(n1705) );
  MXI2X1 U1626 ( .A(n1709), .B(n1710), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_16_), .Y(n7334) );
  AOI21X1 U1627 ( .A0(n1711), .A1(n38), .B0(n75), .Y(n1710) );
  CLKNAND2X2 U1628 ( .A(n25), .B(n1712), .Y(n1709) );
  MXI2X1 U1629 ( .A(n1713), .B(n1714), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_15_), .Y(n7333) );
  AOI2B1X1 U1630 ( .A1N(n1715), .A0(n33), .B0(n82), .Y(n1714) );
  CLKNAND2X2 U1631 ( .A(n25), .B(n1715), .Y(n1713) );
  MXI2X1 U1632 ( .A(n1716), .B(n1717), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_14_), .Y(n7332) );
  AOI21X1 U1633 ( .A0(n1718), .A1(n39), .B0(n74), .Y(n1717) );
  CLKNAND2X2 U1634 ( .A(n24), .B(n1719), .Y(n1716) );
  MXI2X1 U1635 ( .A(n1720), .B(n1721), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_13_), .Y(n7331) );
  AOI21X1 U1636 ( .A0(n1722), .A1(n39), .B0(n74), .Y(n1721) );
  CLKNAND2X2 U1637 ( .A(n24), .B(n1723), .Y(n1720) );
  MXI2X1 U1638 ( .A(n1724), .B(n1725), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_12_), .Y(n7330) );
  AOI21X1 U1639 ( .A0(n1726), .A1(n39), .B0(n74), .Y(n1725) );
  CLKNAND2X2 U1640 ( .A(n24), .B(n1727), .Y(n1724) );
  MXI2X1 U1641 ( .A(n1728), .B(n1729), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_11_), .Y(n7329) );
  AOI21X1 U1642 ( .A0(n1730), .A1(n39), .B0(n74), .Y(n1729) );
  CLKNAND2X2 U1643 ( .A(n24), .B(n1731), .Y(n1728) );
  MXI2X1 U1644 ( .A(n1732), .B(n1733), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_10_), .Y(n7328) );
  AOI21X1 U1645 ( .A0(n1734), .A1(n39), .B0(n74), .Y(n1733) );
  CLKNAND2X2 U1646 ( .A(n24), .B(n1735), .Y(n1732) );
  MXI2X1 U1647 ( .A(n1736), .B(n1737), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_9_), .Y(n7327) );
  AOI21X1 U1648 ( .A0(n1738), .A1(n39), .B0(n74), .Y(n1737) );
  CLKNAND2X2 U1649 ( .A(n24), .B(n1739), .Y(n1736) );
  MXI2X1 U1650 ( .A(n1740), .B(n1741), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_8_), .Y(n7326) );
  AOI21X1 U1651 ( .A0(n1742), .A1(n39), .B0(n74), .Y(n1741) );
  CLKNAND2X2 U1652 ( .A(n24), .B(n1743), .Y(n1740) );
  MXI2X1 U1653 ( .A(n1744), .B(n1745), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_7_), .Y(n7325) );
  AOI21X1 U1654 ( .A0(n1746), .A1(n39), .B0(n74), .Y(n1745) );
  CLKNAND2X2 U1655 ( .A(n23), .B(n1747), .Y(n1744) );
  MXI2X1 U1656 ( .A(n1748), .B(n1749), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_6_), .Y(n7324) );
  AOI21X1 U1657 ( .A0(n1750), .A1(n39), .B0(n74), .Y(n1749) );
  NAND2BX1 U1658 ( .AN(n1750), .B(n35), .Y(n1748) );
  MXI2X1 U1659 ( .A(n1751), .B(n1752), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_5_), .Y(n7323) );
  AOI21X1 U1660 ( .A0(n1753), .A1(n40), .B0(n74), .Y(n1752) );
  NAND2BX1 U1661 ( .AN(n1753), .B(n34), .Y(n1751) );
  MXI2X1 U1662 ( .A(n1754), .B(n1755), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_4_), .Y(n7322) );
  AOI21X1 U1663 ( .A0(n1756), .A1(n40), .B0(n74), .Y(n1755) );
  NAND2BX1 U1664 ( .AN(n1756), .B(n34), .Y(n1754) );
  MXI2X1 U1665 ( .A(n1757), .B(n1758), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_3_), .Y(n7321) );
  AOI21X1 U1666 ( .A0(n1759), .A1(n40), .B0(n74), .Y(n1758) );
  NAND2BX1 U1667 ( .AN(n1759), .B(n34), .Y(n1757) );
  MXI2X1 U1668 ( .A(n1760), .B(n1761), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_2_), .Y(n7320) );
  AOI21X1 U1669 ( .A0(n1762), .A1(n40), .B0(n74), .Y(n1761) );
  NAND2BX1 U1670 ( .AN(n1762), .B(n34), .Y(n1760) );
  MXI2X1 U1671 ( .A(n1763), .B(n1764), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_1_), .Y(n7319) );
  AOI21X1 U1672 ( .A0(n1765), .A1(n40), .B0(n73), .Y(n1764) );
  NAND2BX1 U1673 ( .AN(n1765), .B(n34), .Y(n1763) );
  MXI2X1 U1674 ( .A(n1766), .B(n1767), .S0(
        Inst_forkAE_MainPart1_Tag_Reg_Output_0_), .Y(n7318) );
  AOI21X1 U1675 ( .A0(n1768), .A1(n41), .B0(n73), .Y(n1767) );
  NAND2BX1 U1676 ( .AN(n1768), .B(n34), .Y(n1766) );
  NOR2X1 U1677 ( .A(n82), .B(rst), .Y(n587) );
  AOI211X1 U1678 ( .A0(dec), .A1(done), .B0(n1769), .C0(rst), .Y(n588) );
  CLKINVX1 U1679 ( .A(n1770), .Y(n1769) );
  OAI2B2X1 U1680 ( .A1N(Tag1[127]), .A0(n102), .B0(n1771), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n387) );
  CLKINVX1 U1681 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[127]), .Y(n1771)
         );
  XNOR2X1 U1682 ( .A(n1772), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[127]), 
        .Y(Tag1[127]) );
  OAI2B2X1 U1683 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[126]), .A0(n124), 
        .B0(n566), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n386) );
  XOR2X1 U1684 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[126]), .B(n1773), 
        .Y(n566) );
  OAI2B2X1 U1685 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[125]), .A0(n124), 
        .B0(n567), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n385) );
  XOR2X1 U1686 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[125]), .B(n1774), 
        .Y(n567) );
  OAI2B2X1 U1687 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[124]), .A0(n124), 
        .B0(n568), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n384) );
  XOR2X1 U1688 ( .A(n1775), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[124]), 
        .Y(n568) );
  OAI2B2X1 U1689 ( .A1N(Tag1[123]), .A0(n102), .B0(n1776), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n383) );
  CLKINVX1 U1690 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[123]), .Y(n1776)
         );
  XOR2X1 U1691 ( .A(n1777), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[123]), 
        .Y(Tag1[123]) );
  OAI2B2X1 U1692 ( .A1N(Tag1[122]), .A0(n102), .B0(n1778), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n382) );
  CLKINVX1 U1693 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[122]), .Y(n1778)
         );
  XOR2X1 U1694 ( .A(n1779), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[122]), 
        .Y(Tag1[122]) );
  OAI2B2X1 U1695 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[121]), .A0(n124), 
        .B0(n569), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n381) );
  XOR2X1 U1696 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[121]), .B(n1780), 
        .Y(n569) );
  OAI2B2X1 U1697 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[120]), .A0(n124), 
        .B0(n570), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n380) );
  XOR2X1 U1698 ( .A(n1781), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[120]), 
        .Y(n570) );
  OAI2B2X1 U1699 ( .A1N(Tag1[119]), .A0(n102), .B0(n1782), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n379) );
  CLKINVX1 U1700 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[119]), .Y(n1782)
         );
  XOR2X1 U1701 ( .A(n1783), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[119]), 
        .Y(Tag1[119]) );
  OAI2B2X1 U1702 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[118]), .A0(n124), 
        .B0(n571), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n378) );
  XOR2X1 U1703 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[118]), .B(n1784), 
        .Y(n571) );
  OAI2B2X1 U1704 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[117]), .A0(n124), 
        .B0(n572), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n377) );
  XOR2X1 U1705 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[117]), .B(n1785), 
        .Y(n572) );
  OAI2B2X1 U1706 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[116]), .A0(n124), 
        .B0(n573), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n376) );
  XOR2X1 U1707 ( .A(n1786), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[116]), 
        .Y(n573) );
  OAI2B2X1 U1708 ( .A1N(Tag1[115]), .A0(n102), .B0(n1787), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n375) );
  CLKINVX1 U1709 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[115]), .Y(n1787)
         );
  XOR2X1 U1710 ( .A(n1788), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[115]), 
        .Y(Tag1[115]) );
  OAI2B2X1 U1711 ( .A1N(Tag1[114]), .A0(n103), .B0(n1789), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n374) );
  CLKINVX1 U1712 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[114]), .Y(n1789)
         );
  XOR2X1 U1713 ( .A(n1790), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[114]), 
        .Y(Tag1[114]) );
  OAI2B2X1 U1714 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[113]), .A0(n124), 
        .B0(n574), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n373) );
  XOR2X1 U1715 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[113]), .B(n1791), 
        .Y(n574) );
  OAI2B2X1 U1716 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[112]), .A0(n124), 
        .B0(n575), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n372) );
  XOR2X1 U1717 ( .A(n1792), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[112]), 
        .Y(n575) );
  OAI2B2X1 U1718 ( .A1N(Tag1[111]), .A0(n103), .B0(n1793), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n371) );
  CLKINVX1 U1719 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[111]), .Y(n1793)
         );
  XOR2X1 U1720 ( .A(n1794), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[111]), 
        .Y(Tag1[111]) );
  OAI2B2X1 U1721 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[110]), .A0(n124), 
        .B0(n576), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n370) );
  XOR2X1 U1722 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[110]), .B(n1795), 
        .Y(n576) );
  OAI2B2X1 U1723 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[109]), .A0(n124), 
        .B0(n577), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n369) );
  XOR2X1 U1724 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[109]), .B(n1796), 
        .Y(n577) );
  OAI2B2X1 U1725 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[108]), .A0(n124), 
        .B0(n578), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n368) );
  XOR2X1 U1726 ( .A(n1797), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[108]), 
        .Y(n578) );
  OAI2B2X1 U1727 ( .A1N(Tag1[107]), .A0(n103), .B0(n1798), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n367) );
  CLKINVX1 U1728 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[107]), .Y(n1798)
         );
  XOR2X1 U1729 ( .A(n1799), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[107]), 
        .Y(Tag1[107]) );
  OAI2B2X1 U1730 ( .A1N(Tag1[106]), .A0(n103), .B0(n1800), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n366) );
  CLKINVX1 U1731 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[106]), .Y(n1800)
         );
  XOR2X1 U1732 ( .A(n1801), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[106]), 
        .Y(Tag1[106]) );
  OAI2B2X1 U1733 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[105]), .A0(n125), 
        .B0(n579), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n365) );
  XOR2X1 U1734 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[105]), .B(n1802), 
        .Y(n579) );
  OAI2B2X1 U1735 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[104]), .A0(n125), 
        .B0(n580), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n364) );
  XOR2X1 U1736 ( .A(n1803), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[104]), 
        .Y(n580) );
  OAI2B2X1 U1737 ( .A1N(Tag1[103]), .A0(n103), .B0(n1804), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n363) );
  CLKINVX1 U1738 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[103]), .Y(n1804)
         );
  XOR2X1 U1739 ( .A(n1805), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[103]), 
        .Y(Tag1[103]) );
  OAI2B2X1 U1740 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[102]), .A0(n125), 
        .B0(n581), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n362) );
  XOR2X1 U1741 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[102]), .B(n1806), 
        .Y(n581) );
  OAI2B2X1 U1742 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[101]), .A0(n125), 
        .B0(n582), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n361) );
  XOR2X1 U1743 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[101]), .B(n1807), 
        .Y(n582) );
  OAI2B2X1 U1744 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[100]), .A0(n125), 
        .B0(n583), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n360) );
  XOR2X1 U1745 ( .A(n1808), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[100]), 
        .Y(n583) );
  OAI2B2X1 U1746 ( .A1N(Tag1[99]), .A0(n103), .B0(n1809), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n359) );
  CLKINVX1 U1747 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[99]), .Y(n1809) );
  XOR2X1 U1748 ( .A(n1810), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[99]), .Y(
        Tag1[99]) );
  OAI2B2X1 U1749 ( .A1N(Tag1[98]), .A0(n103), .B0(n1811), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n358) );
  CLKINVX1 U1750 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[98]), .Y(n1811) );
  XOR2X1 U1751 ( .A(n1812), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[98]), .Y(
        Tag1[98]) );
  OAI2B2X1 U1752 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[97]), .A0(n125), 
        .B0(n528), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n357) );
  XOR2X1 U1753 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[97]), .B(n1813), .Y(
        n528) );
  OAI2B2X1 U1754 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[96]), .A0(n125), 
        .B0(n529), .B1(n108), .Y(Inst_forkAE_MainPart1_AuthRegInst_n356) );
  XOR2X1 U1755 ( .A(n1814), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[96]), .Y(
        n529) );
  OAI2B2X1 U1756 ( .A1N(Tag1[95]), .A0(n107), .B0(n1815), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n355) );
  CLKINVX1 U1757 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[95]), .Y(n1815) );
  XOR2X1 U1758 ( .A(n1816), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[95]), .Y(
        Tag1[95]) );
  OAI2B2X1 U1759 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[94]), .A0(n125), 
        .B0(n530), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n354) );
  XOR2X1 U1760 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[94]), .B(n1817), .Y(
        n530) );
  OAI2B2X1 U1761 ( .A1N(Tag1[93]), .A0(n107), .B0(n1818), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n353) );
  CLKINVX1 U1762 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[93]), .Y(n1818) );
  XOR2X1 U1763 ( .A(n1819), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[93]), .Y(
        Tag1[93]) );
  OAI2B2X1 U1764 ( .A1N(Tag1[92]), .A0(n107), .B0(n1820), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n352) );
  CLKINVX1 U1765 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[92]), .Y(n1820) );
  XNOR2X1 U1766 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[92]), .B(n1821), 
        .Y(Tag1[92]) );
  OAI2B2X1 U1767 ( .A1N(Tag1[91]), .A0(n107), .B0(n1822), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n351) );
  CLKINVX1 U1768 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[91]), .Y(n1822) );
  XOR2X1 U1769 ( .A(n1823), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[91]), .Y(
        Tag1[91]) );
  OAI2B2X1 U1770 ( .A1N(Tag1[90]), .A0(n107), .B0(n1824), .B1(n134), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n350) );
  CLKINVX1 U1771 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[90]), .Y(n1824) );
  XOR2X1 U1772 ( .A(n1825), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[90]), .Y(
        Tag1[90]) );
  OAI2B2X1 U1773 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[89]), .A0(n125), 
        .B0(n531), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n349) );
  XOR2X1 U1774 ( .A(n1826), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[89]), .Y(
        n531) );
  OAI2B2X1 U1775 ( .A1N(Tag1[88]), .A0(n108), .B0(n1827), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n348) );
  CLKINVX1 U1776 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[88]), .Y(n1827) );
  XNOR2X1 U1777 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[88]), .B(n1828), 
        .Y(Tag1[88]) );
  OAI2B2X1 U1778 ( .A1N(Tag1[87]), .A0(n107), .B0(n1829), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n347) );
  CLKINVX1 U1779 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[87]), .Y(n1829) );
  XOR2X1 U1780 ( .A(n1830), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[87]), .Y(
        Tag1[87]) );
  OAI2B2X1 U1781 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[86]), .A0(n125), 
        .B0(n532), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n346) );
  XOR2X1 U1782 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[86]), .B(n1831), .Y(
        n532) );
  OAI2B2X1 U1783 ( .A1N(Tag1[85]), .A0(n108), .B0(n1832), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n345) );
  CLKINVX1 U1784 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[85]), .Y(n1832) );
  XOR2X1 U1785 ( .A(n1833), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[85]), .Y(
        Tag1[85]) );
  OAI2B2X1 U1786 ( .A1N(Tag1[84]), .A0(n107), .B0(n1834), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n344) );
  CLKINVX1 U1787 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[84]), .Y(n1834) );
  XNOR2X1 U1788 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[84]), .B(n1835), 
        .Y(Tag1[84]) );
  OAI2B2X1 U1789 ( .A1N(Tag1[83]), .A0(n107), .B0(n1836), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n343) );
  CLKINVX1 U1790 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[83]), .Y(n1836) );
  XOR2X1 U1791 ( .A(n1837), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[83]), .Y(
        Tag1[83]) );
  OAI2B2X1 U1792 ( .A1N(Tag1[82]), .A0(n107), .B0(n1838), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n342) );
  CLKINVX1 U1793 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[82]), .Y(n1838) );
  XOR2X1 U1794 ( .A(n1839), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[82]), .Y(
        Tag1[82]) );
  OAI2B2X1 U1795 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[81]), .A0(n125), 
        .B0(n533), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n341) );
  XOR2X1 U1796 ( .A(n1840), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[81]), .Y(
        n533) );
  OAI2B2X1 U1797 ( .A1N(Tag1[80]), .A0(n107), .B0(n1841), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n340) );
  CLKINVX1 U1798 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[80]), .Y(n1841) );
  XNOR2X1 U1799 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[80]), .B(n1842), 
        .Y(Tag1[80]) );
  OAI2B2X1 U1800 ( .A1N(Tag1[79]), .A0(n107), .B0(n1843), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n339) );
  CLKINVX1 U1801 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[79]), .Y(n1843) );
  XOR2X1 U1802 ( .A(n1844), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[79]), .Y(
        Tag1[79]) );
  OAI2B2X1 U1803 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[78]), .A0(n125), 
        .B0(n534), .B1(n115), .Y(Inst_forkAE_MainPart1_AuthRegInst_n338) );
  XOR2X1 U1804 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[78]), .B(n1845), .Y(
        n534) );
  OAI2B2X1 U1805 ( .A1N(Tag1[77]), .A0(n107), .B0(n1846), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n337) );
  CLKINVX1 U1806 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[77]), .Y(n1846) );
  XOR2X1 U1807 ( .A(n1847), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[77]), .Y(
        Tag1[77]) );
  OAI2B2X1 U1808 ( .A1N(Tag1[76]), .A0(n107), .B0(n1848), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n336) );
  CLKINVX1 U1809 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[76]), .Y(n1848) );
  XNOR2X1 U1810 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[76]), .B(n1849), 
        .Y(Tag1[76]) );
  OAI2B2X1 U1811 ( .A1N(Tag1[75]), .A0(n106), .B0(n1850), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n335) );
  CLKINVX1 U1812 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[75]), .Y(n1850) );
  XOR2X1 U1813 ( .A(n1851), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[75]), .Y(
        Tag1[75]) );
  OAI2B2X1 U1814 ( .A1N(Tag1[74]), .A0(n106), .B0(n1852), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n334) );
  CLKINVX1 U1815 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[74]), .Y(n1852) );
  XOR2X1 U1816 ( .A(n1853), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[74]), .Y(
        Tag1[74]) );
  OAI2B2X1 U1817 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[73]), .A0(n126), 
        .B0(n535), .B1(n115), .Y(Inst_forkAE_MainPart1_AuthRegInst_n333) );
  XOR2X1 U1818 ( .A(n1854), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[73]), .Y(
        n535) );
  OAI2B2X1 U1819 ( .A1N(Tag1[72]), .A0(n106), .B0(n1855), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n332) );
  CLKINVX1 U1820 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[72]), .Y(n1855) );
  XNOR2X1 U1821 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[72]), .B(n1856), 
        .Y(Tag1[72]) );
  OAI2B2X1 U1822 ( .A1N(Tag1[71]), .A0(n106), .B0(n1857), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n331) );
  CLKINVX1 U1823 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[71]), .Y(n1857) );
  XOR2X1 U1824 ( .A(n1858), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[71]), .Y(
        Tag1[71]) );
  OAI2B2X1 U1825 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[70]), .A0(n126), 
        .B0(n536), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n330) );
  XOR2X1 U1826 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[70]), .B(n1859), .Y(
        n536) );
  OAI2B2X1 U1827 ( .A1N(Tag1[69]), .A0(n106), .B0(n1860), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n329) );
  CLKINVX1 U1828 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[69]), .Y(n1860) );
  XOR2X1 U1829 ( .A(n1861), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[69]), .Y(
        Tag1[69]) );
  OAI2B2X1 U1830 ( .A1N(Tag1[68]), .A0(n106), .B0(n1862), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n328) );
  CLKINVX1 U1831 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[68]), .Y(n1862) );
  XNOR2X1 U1832 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[68]), .B(n1863), 
        .Y(Tag1[68]) );
  OAI2B2X1 U1833 ( .A1N(Tag1[67]), .A0(n106), .B0(n1864), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n327) );
  CLKINVX1 U1834 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[67]), .Y(n1864) );
  XOR2X1 U1835 ( .A(n1865), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[67]), .Y(
        Tag1[67]) );
  OAI2B2X1 U1836 ( .A1N(Tag1[66]), .A0(n106), .B0(n1866), .B1(n135), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n326) );
  CLKINVX1 U1837 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[66]), .Y(n1866) );
  XOR2X1 U1838 ( .A(n1867), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[66]), .Y(
        Tag1[66]) );
  OAI2B2X1 U1839 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[65]), .A0(n126), 
        .B0(n538), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n325) );
  XOR2X1 U1840 ( .A(n1868), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[65]), .Y(
        n538) );
  OAI2B2X1 U1841 ( .A1N(Tag1[64]), .A0(n106), .B0(n1869), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n324) );
  CLKINVX1 U1842 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[64]), .Y(n1869) );
  XNOR2X1 U1843 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[64]), .B(n1870), 
        .Y(Tag1[64]) );
  OAI2B2X1 U1844 ( .A1N(Tag1[63]), .A0(n106), .B0(n1871), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n323) );
  CLKINVX1 U1845 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[63]), .Y(n1871) );
  XOR2X1 U1846 ( .A(n1872), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[63]), .Y(
        Tag1[63]) );
  OAI2B2X1 U1847 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[62]), .A0(n126), 
        .B0(n539), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n322) );
  XOR2X1 U1848 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[62]), .B(n1873), .Y(
        n539) );
  OAI2B2X1 U1849 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[61]), .A0(n126), 
        .B0(n540), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n321) );
  XOR2X1 U1850 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[61]), .B(n1874), .Y(
        n540) );
  OAI2B2X1 U1851 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[60]), .A0(n126), 
        .B0(n541), .B1(n114), .Y(Inst_forkAE_MainPart1_AuthRegInst_n320) );
  XOR2X1 U1852 ( .A(n1875), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[60]), .Y(
        n541) );
  OAI2B2X1 U1853 ( .A1N(Tag1[59]), .A0(n106), .B0(n1876), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n319) );
  CLKINVX1 U1854 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[59]), .Y(n1876) );
  XOR2X1 U1855 ( .A(n1877), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[59]), .Y(
        Tag1[59]) );
  OAI2B2X1 U1856 ( .A1N(Tag1[58]), .A0(n106), .B0(n1878), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n318) );
  CLKINVX1 U1857 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[58]), .Y(n1878) );
  XOR2X1 U1858 ( .A(n1879), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[58]), .Y(
        Tag1[58]) );
  OAI2B2X1 U1859 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[57]), .A0(n128), 
        .B0(n542), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n317) );
  XOR2X1 U1860 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[57]), .B(n1880), .Y(
        n542) );
  OAI2B2X1 U1861 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[56]), .A0(n129), 
        .B0(n543), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n316) );
  XOR2X1 U1862 ( .A(n1881), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[56]), .Y(
        n543) );
  OAI2B2X1 U1863 ( .A1N(Tag1[55]), .A0(n105), .B0(n1882), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n315) );
  CLKINVX1 U1864 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[55]), .Y(n1882) );
  XOR2X1 U1865 ( .A(n1883), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[55]), .Y(
        Tag1[55]) );
  OAI2B2X1 U1866 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[54]), .A0(n128), 
        .B0(n544), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n314) );
  XOR2X1 U1867 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[54]), .B(n1884), .Y(
        n544) );
  OAI2B2X1 U1868 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[53]), .A0(n129), 
        .B0(n545), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n313) );
  XOR2X1 U1869 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[53]), .B(n1885), .Y(
        n545) );
  OAI2B2X1 U1870 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[52]), .A0(n128), 
        .B0(n546), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n312) );
  XOR2X1 U1871 ( .A(n1886), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[52]), .Y(
        n546) );
  OAI2B2X1 U1872 ( .A1N(Tag1[51]), .A0(n105), .B0(n1887), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n311) );
  CLKINVX1 U1873 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[51]), .Y(n1887) );
  XOR2X1 U1874 ( .A(n1888), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[51]), .Y(
        Tag1[51]) );
  OAI2B2X1 U1875 ( .A1N(Tag1[50]), .A0(n105), .B0(n1889), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n310) );
  CLKINVX1 U1876 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[50]), .Y(n1889) );
  XOR2X1 U1877 ( .A(n1890), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[50]), .Y(
        Tag1[50]) );
  OAI2B2X1 U1878 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[49]), .A0(n128), 
        .B0(n547), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n309) );
  XOR2X1 U1879 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[49]), .B(n1891), .Y(
        n547) );
  OAI2B2X1 U1880 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[48]), .A0(n128), 
        .B0(n548), .B1(n113), .Y(Inst_forkAE_MainPart1_AuthRegInst_n308) );
  XOR2X1 U1881 ( .A(n1892), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[48]), .Y(
        n548) );
  OAI2B2X1 U1882 ( .A1N(Tag1[47]), .A0(n105), .B0(n1893), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n307) );
  CLKINVX1 U1883 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[47]), .Y(n1893) );
  XOR2X1 U1884 ( .A(n1894), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[47]), .Y(
        Tag1[47]) );
  OAI2B2X1 U1885 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[46]), .A0(n128), 
        .B0(n549), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n306) );
  XOR2X1 U1886 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[46]), .B(n1895), .Y(
        n549) );
  OAI2B2X1 U1887 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[45]), .A0(n128), 
        .B0(n550), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n305) );
  XOR2X1 U1888 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[45]), .B(n1896), .Y(
        n550) );
  OAI2B2X1 U1889 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[44]), .A0(n128), 
        .B0(n551), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n304) );
  XOR2X1 U1890 ( .A(n1897), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[44]), .Y(
        n551) );
  OAI2B2X1 U1891 ( .A1N(Tag1[43]), .A0(n105), .B0(n1898), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n303) );
  CLKINVX1 U1892 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[43]), .Y(n1898) );
  XOR2X1 U1893 ( .A(n1899), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[43]), .Y(
        Tag1[43]) );
  OAI2B2X1 U1894 ( .A1N(Tag1[42]), .A0(n105), .B0(n1900), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n302) );
  CLKINVX1 U1895 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[42]), .Y(n1900) );
  XOR2X1 U1896 ( .A(n1901), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[42]), .Y(
        Tag1[42]) );
  OAI2B2X1 U1897 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[41]), .A0(n128), 
        .B0(n552), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n301) );
  XOR2X1 U1898 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[41]), .B(n1902), .Y(
        n552) );
  OAI2B2X1 U1899 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[40]), .A0(n128), 
        .B0(n553), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n300) );
  XOR2X1 U1900 ( .A(n1903), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[40]), .Y(
        n553) );
  OAI2B2X1 U1901 ( .A1N(Tag1[39]), .A0(n105), .B0(n1904), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n299) );
  CLKINVX1 U1902 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[39]), .Y(n1904) );
  XOR2X1 U1903 ( .A(n1905), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[39]), .Y(
        Tag1[39]) );
  OAI2B2X1 U1904 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[38]), .A0(n128), 
        .B0(n554), .B1(n112), .Y(Inst_forkAE_MainPart1_AuthRegInst_n298) );
  XOR2X1 U1905 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[38]), .B(n1906), .Y(
        n554) );
  OAI2B2X1 U1906 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[37]), .A0(n128), 
        .B0(n555), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n297) );
  XOR2X1 U1907 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[37]), .B(n1907), .Y(
        n555) );
  OAI2B2X1 U1908 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[36]), .A0(n127), 
        .B0(n556), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n296) );
  XOR2X1 U1909 ( .A(n1908), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[36]), .Y(
        n556) );
  OAI2B2X1 U1910 ( .A1N(Tag1[35]), .A0(n105), .B0(n1909), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n295) );
  CLKINVX1 U1911 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[35]), .Y(n1909) );
  XOR2X1 U1912 ( .A(n1910), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[35]), .Y(
        Tag1[35]) );
  OAI2B2X1 U1913 ( .A1N(Tag1[34]), .A0(n105), .B0(n1911), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n294) );
  CLKINVX1 U1914 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[34]), .Y(n1911) );
  XOR2X1 U1915 ( .A(n1912), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[34]), .Y(
        Tag1[34]) );
  OAI2B2X1 U1916 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[33]), .A0(n127), 
        .B0(n557), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n293) );
  XOR2X1 U1917 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[33]), .B(n1913), .Y(
        n557) );
  OAI2B2X1 U1918 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[32]), .A0(n127), 
        .B0(n558), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n292) );
  XOR2X1 U1919 ( .A(n1914), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[32]), .Y(
        n558) );
  OAI2B2X1 U1920 ( .A1N(Tag1[31]), .A0(n105), .B0(n1915), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n291) );
  CLKINVX1 U1921 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[31]), .Y(n1915) );
  XOR2X1 U1922 ( .A(n1916), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[31]), .Y(
        Tag1[31]) );
  OAI2B2X1 U1923 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[30]), .A0(n127), 
        .B0(n559), .B1(n111), .Y(Inst_forkAE_MainPart1_AuthRegInst_n290) );
  XOR2X1 U1924 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[30]), .B(n1917), .Y(
        n559) );
  OAI2B2X1 U1925 ( .A1N(Tag1[29]), .A0(n105), .B0(n1918), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n289) );
  CLKINVX1 U1926 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[29]), .Y(n1918) );
  XOR2X1 U1927 ( .A(n1919), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[29]), .Y(
        Tag1[29]) );
  OAI2B2X1 U1928 ( .A1N(Tag1[28]), .A0(n105), .B0(n1920), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n288) );
  CLKINVX1 U1929 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[28]), .Y(n1920) );
  XNOR2X1 U1930 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[28]), .B(n1921), 
        .Y(Tag1[28]) );
  OAI2B2X1 U1931 ( .A1N(Tag1[27]), .A0(n105), .B0(n1922), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n287) );
  CLKINVX1 U1932 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[27]), .Y(n1922) );
  XOR2X1 U1933 ( .A(n1923), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[27]), .Y(
        Tag1[27]) );
  OAI2B2X1 U1934 ( .A1N(Tag1[26]), .A0(n104), .B0(n1924), .B1(n136), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n286) );
  CLKINVX1 U1935 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[26]), .Y(n1924) );
  XOR2X1 U1936 ( .A(n1925), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[26]), .Y(
        Tag1[26]) );
  OAI2B2X1 U1937 ( .A1N(Tag1[25]), .A0(n104), .B0(n1926), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n285) );
  CLKINVX1 U1938 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[25]), .Y(n1926) );
  XNOR2X1 U1939 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[25]), .B(n1927), 
        .Y(Tag1[25]) );
  OAI2B2X1 U1940 ( .A1N(Tag1[24]), .A0(n104), .B0(n1928), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n284) );
  CLKINVX1 U1941 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[24]), .Y(n1928) );
  XNOR2X1 U1942 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[24]), .B(n1929), 
        .Y(Tag1[24]) );
  OAI2B2X1 U1943 ( .A1N(Tag1[23]), .A0(n106), .B0(n1930), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n283) );
  CLKINVX1 U1944 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[23]), .Y(n1930) );
  XOR2X1 U1945 ( .A(n1931), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[23]), .Y(
        Tag1[23]) );
  OAI2B2X1 U1946 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[22]), .A0(n127), 
        .B0(n560), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n282) );
  XOR2X1 U1947 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[22]), .B(n1932), .Y(
        n560) );
  OAI2B2X1 U1948 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[21]), .A0(n127), 
        .B0(n561), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n281) );
  XOR2X1 U1949 ( .A(n1933), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[21]), .Y(
        n561) );
  OAI2B2X1 U1950 ( .A1N(Tag1[20]), .A0(n104), .B0(n1934), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n280) );
  CLKINVX1 U1951 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[20]), .Y(n1934) );
  XNOR2X1 U1952 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[20]), .B(n1935), 
        .Y(Tag1[20]) );
  OAI2B2X1 U1953 ( .A1N(Tag1[19]), .A0(n104), .B0(n1936), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n279) );
  CLKINVX1 U1954 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[19]), .Y(n1936) );
  XOR2X1 U1955 ( .A(n1937), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[19]), .Y(
        Tag1[19]) );
  OAI2B2X1 U1956 ( .A1N(Tag1[18]), .A0(n104), .B0(n1938), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n278) );
  CLKINVX1 U1957 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[18]), .Y(n1938) );
  XOR2X1 U1958 ( .A(n1939), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[18]), .Y(
        Tag1[18]) );
  OAI2B2X1 U1959 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[17]), .A0(n127), 
        .B0(n563), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n277) );
  XOR2X1 U1960 ( .A(n1940), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[17]), .Y(
        n563) );
  OAI2B2X1 U1961 ( .A1N(Tag1[16]), .A0(n104), .B0(n1941), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n276) );
  CLKINVX1 U1962 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[16]), .Y(n1941) );
  XNOR2X1 U1963 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[16]), .B(n1942), 
        .Y(Tag1[16]) );
  OAI2B2X1 U1964 ( .A1N(Tag1[15]), .A0(n104), .B0(n1943), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n275) );
  CLKINVX1 U1965 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[15]), .Y(n1943) );
  XOR2X1 U1966 ( .A(n1944), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[15]), .Y(
        Tag1[15]) );
  OAI2B2X1 U1967 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[14]), .A0(n127), 
        .B0(n564), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n274) );
  XOR2X1 U1968 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[14]), .B(n1945), .Y(
        n564) );
  OAI2B2X1 U1969 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[13]), .A0(n127), 
        .B0(n565), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n273) );
  XOR2X1 U1970 ( .A(n1946), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[13]), .Y(
        n565) );
  OAI2B2X1 U1971 ( .A1N(Tag1[12]), .A0(n104), .B0(n1947), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n272) );
  CLKINVX1 U1972 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[12]), .Y(n1947) );
  XNOR2X1 U1973 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[12]), .B(n1948), 
        .Y(Tag1[12]) );
  OAI2B2X1 U1974 ( .A1N(Tag1[11]), .A0(n104), .B0(n1949), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n271) );
  CLKINVX1 U1975 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[11]), .Y(n1949) );
  XOR2X1 U1976 ( .A(n1950), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[11]), .Y(
        Tag1[11]) );
  OAI2B2X1 U1977 ( .A1N(Tag1[10]), .A0(n104), .B0(n1951), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n270) );
  CLKINVX1 U1978 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[10]), .Y(n1951) );
  XOR2X1 U1979 ( .A(n1952), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[10]), .Y(
        Tag1[10]) );
  OAI2B2X1 U1980 ( .A1N(Tag1[9]), .A0(n104), .B0(n1953), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n269) );
  CLKINVX1 U1981 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[9]), .Y(n1953) );
  XNOR2X1 U1982 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[9]), .B(n1954), .Y(
        Tag1[9]) );
  OAI2B2X1 U1983 ( .A1N(Tag1[8]), .A0(n104), .B0(n1955), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n268) );
  CLKINVX1 U1984 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[8]), .Y(n1955) );
  XNOR2X1 U1985 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[8]), .B(n1956), .Y(
        Tag1[8]) );
  OAI2B2X1 U1986 ( .A1N(Tag1[7]), .A0(n103), .B0(n1957), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n267) );
  CLKINVX1 U1987 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[7]), .Y(n1957) );
  XOR2X1 U1988 ( .A(n1958), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[7]), .Y(
        Tag1[7]) );
  OAI2B2X1 U1989 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[6]), .A0(n126), 
        .B0(n537), .B1(n109), .Y(Inst_forkAE_MainPart1_AuthRegInst_n266) );
  XOR2X1 U1990 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[6]), .B(n1959), .Y(
        n537) );
  OAI2B2X1 U1991 ( .A1N(Tag1[5]), .A0(n103), .B0(n1960), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n265) );
  CLKINVX1 U1992 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[5]), .Y(n1960) );
  XOR2X1 U1993 ( .A(n1961), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[5]), .Y(
        Tag1[5]) );
  OAI2B2X1 U1994 ( .A1N(Tag1[4]), .A0(n103), .B0(n1962), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n264) );
  CLKINVX1 U1995 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[4]), .Y(n1962) );
  XNOR2X1 U1996 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[4]), .B(n1963), .Y(
        Tag1[4]) );
  OAI2B2X1 U1997 ( .A1N(Tag1[3]), .A0(n103), .B0(n1964), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n263) );
  CLKINVX1 U1998 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[3]), .Y(n1964) );
  XOR2X1 U1999 ( .A(n1965), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[3]), .Y(
        Tag1[3]) );
  OAI2B2X1 U2000 ( .A1N(Tag1[2]), .A0(n103), .B0(n1966), .B1(n137), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n262) );
  CLKINVX1 U2001 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[2]), .Y(n1966) );
  XOR2X1 U2002 ( .A(n1967), .B(Inst_forkAE_MainPart1_Auth_Reg_Output[2]), .Y(
        Tag1[2]) );
  OAI2B2X1 U2003 ( .A1N(Inst_forkAE_MainPart1_Auth_Reg_Output[1]), .A0(n126), 
        .B0(n562), .B1(n110), .Y(Inst_forkAE_MainPart1_AuthRegInst_n261) );
  XOR2X1 U2004 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[1]), .B(n1968), .Y(
        n562) );
  OAI2B2X1 U2005 ( .A1N(Tag1[0]), .A0(n96), .B0(n1969), .B1(n131), .Y(
        Inst_forkAE_MainPart1_AuthRegInst_n260) );
  CLKINVX1 U2006 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[0]), .Y(n1969) );
  CLKNAND2X2 U2007 ( .A(n123), .B(n1970), .Y(n1069) );
  OAI21X1 U2008 ( .A0(n1971), .A1(n1972), .B0(n1970), .Y(n1071) );
  XNOR2X1 U2009 ( .A(Inst_forkAE_MainPart1_Auth_Reg_Output[0]), .B(n1973), .Y(
        Tag1[0]) );
  OAI22X1 U2010 ( .A0(Inst_forkAE_LFSRInst_n52), .A1(n1974), .B0(n1975), .B1(
        n1976), .Y(Inst_forkAE_LFSRInst_n63) );
  XOR2X1 U2011 ( .A(n484), .B(Inst_forkAE_CipherInst_TK1_DEC_48_), .Y(n1976)
         );
  OAI22X1 U2012 ( .A0(n1974), .A1(n1977), .B0(n1978), .B1(n1975), .Y(
        Inst_forkAE_LFSRInst_n62) );
  XOR2X1 U2013 ( .A(n465), .B(n3), .Y(n1978) );
  OAI22X1 U2014 ( .A0(Inst_forkAE_LFSRInst_n51), .A1(n1974), .B0(n1975), .B1(
        n1979), .Y(Inst_forkAE_LFSRInst_n61) );
  XOR2X1 U2015 ( .A(n484), .B(Inst_forkAE_CipherInst_TK1_DEC_51_), .Y(n1979)
         );
  CLKNAND2X2 U2016 ( .A(n5715), .B(done), .Y(n1975) );
  CLKINVX1 U2017 ( .A(n1971), .Y(done) );
  CLKNAND2X2 U2018 ( .A(n5715), .B(n1971), .Y(n1974) );
  AOI31X1 U2019 ( .A0(n1980), .A1(n1981), .A2(n1982), .B0(rst), .Y(n5715) );
  CLKINVX1 U2020 ( .A(Inst_forkAE_ControlInst_encdec_started), .Y(n1981) );
  AOI21X1 U2021 ( .A0(n1971), .A1(n1983), .B0(rst), .Y(
        Inst_forkAE_ControlInst_n33) );
  OAI22X1 U2022 ( .A0(a_data), .A1(n1982), .B0(n1980), .B1(n1984), .Y(n1983)
         );
  NOR2X1 U2023 ( .A(n145), .B(n1986), .Y(n1984) );
  CLKNAND2X2 U2024 ( .A(n1987), .B(n1988), .Y(n1971) );
  AOI211X1 U2025 ( .A0(n1989), .A1(Inst_forkAE_CipherInst_ROUND_CST[2]), .B0(
        n1990), .C0(n5718), .Y(n1988) );
  NAND3XL U2026 ( .A(n1991), .B(n1986), .C(n1992), .Y(n1990) );
  NOR4X1 U2027 ( .A(n1993), .B(n1994), .C(n145), .D(n1995), .Y(n1987) );
  MXI2X1 U2028 ( .A(n1989), .B(Inst_forkAE_CipherInst_ROUND_CST[2]), .S0(n1996), .Y(n1995) );
  NOR2X1 U2029 ( .A(rst), .B(n1997), .Y(Inst_forkAE_ControlInst_n32) );
  AOI2BB1X1 U2030 ( .A0N(n159), .A1N(n1998), .B0(n1999), .Y(n1997) );
  AOI21X1 U2031 ( .A0(n2000), .A1(Inst_forkAE_ControlInst_fsm_state_1_), .B0(
        n1986), .Y(n1999) );
  OAI21X1 U2032 ( .A0(rst), .A1(n2001), .B0(n1770), .Y(
        Inst_forkAE_ControlInst_n31) );
  NAND3XL U2033 ( .A(n1980), .B(n1970), .C(enc), .Y(n1770) );
  CLKINVX1 U2034 ( .A(rst), .Y(n1970) );
  AOI21X1 U2035 ( .A0(dec), .A1(n1980), .B0(
        Inst_forkAE_ControlInst_encdec_started), .Y(n2001) );
  NOR2X1 U2036 ( .A(Inst_forkAE_ControlInst_fsm_state_0_), .B(
        Inst_forkAE_ControlInst_fsm_state_1_), .Y(n1980) );
  CLKINVX1 U2037 ( .A(n1992), .Y(Inst_forkAE_CipherInst_ROUND_CST[5]) );
  CLKINVX1 U2038 ( .A(n1991), .Y(Inst_forkAE_CipherInst_ROUND_CST[4]) );
  OAI33X1 U2039 ( .A0(n2002), .A1(n2003), .A2(n2004), .B0(n2005), .B1(n2006), 
        .B2(n2007), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N9) );
  OAI33X1 U2040 ( .A0(n2002), .A1(n2008), .A2(n2009), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .B2(n2010), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N8) );
  OAI33X1 U2041 ( .A0(n2002), .A1(n2011), .A2(n2012), .B0(n2005), .B1(n2013), 
        .B2(n2014), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N7) );
  OAI33X1 U2042 ( .A0(n2002), .A1(n2015), .A2(n2016), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .B2(n2017), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N6) );
  OAI33X1 U2043 ( .A0(n2002), .A1(n2018), .A2(n2019), .B0(n2005), .B1(n2020), 
        .B2(n2021), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N5) );
  OAI33X1 U2044 ( .A0(n2002), .A1(n2022), .A2(n2023), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .B2(n2024), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N4) );
  CLKINVX1 U2045 ( .A(n2025), .Y(n2023) );
  OAI33X1 U2046 ( .A0(n2002), .A1(n2026), .A2(n2027), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .B2(n2028), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N34) );
  CLKINVX1 U2047 ( .A(n2029), .Y(n2027) );
  OAI33X1 U2048 ( .A0(n2002), .A1(n2030), .A2(n2031), .B0(n2005), .B1(n2032), 
        .B2(n2033), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N33) );
  OAI33X1 U2049 ( .A0(n2002), .A1(n2034), .A2(n2035), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .B2(n2036), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N32) );
  CLKINVX1 U2050 ( .A(n2037), .Y(n2035) );
  OAI33X1 U2051 ( .A0(n2002), .A1(n2038), .A2(n2039), .B0(n2005), .B1(n2040), 
        .B2(n2041), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N31) );
  OAI33X1 U2052 ( .A0(n2002), .A1(n2042), .A2(n2043), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .B2(n2044), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N30) );
  CLKINVX1 U2053 ( .A(n2045), .Y(n2043) );
  OAI33X1 U2054 ( .A0(n2002), .A1(n2046), .A2(n2047), .B0(n2005), .B1(n2048), 
        .B2(n2049), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N3) );
  OAI33X1 U2055 ( .A0(n2002), .A1(n2050), .A2(n2051), .B0(n2005), .B1(n2052), 
        .B2(n2053), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N29) );
  OAI33X1 U2056 ( .A0(n2002), .A1(n2054), .A2(n2055), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .B2(n2056), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N28) );
  CLKINVX1 U2057 ( .A(n2057), .Y(n2055) );
  OAI33X1 U2058 ( .A0(n2002), .A1(n2058), .A2(n2059), .B0(n2005), .B1(n2060), 
        .B2(n2061), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N27) );
  OAI33X1 U2059 ( .A0(n2002), .A1(n2062), .A2(n2063), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .B2(n2064), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N26) );
  OAI33X1 U2060 ( .A0(n2002), .A1(n2065), .A2(n2066), .B0(n2005), .B1(n2067), 
        .B2(n2068), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N25) );
  OAI33X1 U2061 ( .A0(n2002), .A1(n2069), .A2(n2070), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .B2(n2071), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N24) );
  OAI33X1 U2062 ( .A0(n2002), .A1(n2072), .A2(n2073), .B0(n2005), .B1(n2074), 
        .B2(n2075), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N23) );
  OAI33X1 U2063 ( .A0(n2002), .A1(n2076), .A2(n2077), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .B2(n2078), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N22) );
  OAI33X1 U2064 ( .A0(n2002), .A1(n2079), .A2(n2080), .B0(n2005), .B1(n2081), 
        .B2(n2082), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N21) );
  OAI33X1 U2065 ( .A0(n2002), .A1(n2083), .A2(n2084), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .B2(n2085), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N20) );
  OAI33X1 U2066 ( .A0(n2002), .A1(n2086), .A2(n2087), .B0(n2005), .B1(n2088), 
        .B2(n2089), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N19) );
  OAI33X1 U2067 ( .A0(n2002), .A1(n2090), .A2(n2091), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .B2(n2092), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N18) );
  OAI33X1 U2068 ( .A0(n2002), .A1(n2093), .A2(n2094), .B0(n2005), .B1(n2095), 
        .B2(n2096), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N17) );
  OAI33X1 U2069 ( .A0(n2002), .A1(n2097), .A2(n2098), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .B2(n2099), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N16) );
  OAI33X1 U2070 ( .A0(n2002), .A1(n2100), .A2(n2101), .B0(n2005), .B1(n2102), 
        .B2(n2103), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N15) );
  OAI33X1 U2071 ( .A0(n2002), .A1(n2104), .A2(n2105), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .B2(n2106), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N14) );
  OAI33X1 U2072 ( .A0(n2002), .A1(n2107), .A2(n2108), .B0(n2005), .B1(n2109), 
        .B2(n2110), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N13) );
  OAI33X1 U2073 ( .A0(n2002), .A1(n2111), .A2(n2112), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .B2(n2113), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N12) );
  OAI33X1 U2074 ( .A0(n2002), .A1(n2114), .A2(n2115), .B0(n2005), .B1(n2116), 
        .B2(n2117), .Y(Inst_forkAE_CipherInst_RF_RS_EX2_N11) );
  OAI33X1 U2075 ( .A0(n2002), .A1(n2118), .A2(n2119), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .B2(n2120), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX2_N10) );
  OAI33X1 U2076 ( .A0(n2002), .A1(n2121), .A2(n2122), .B0(n2005), .B1(n2123), 
        .B2(n2124), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N9) );
  OAI33X1 U2077 ( .A0(n2002), .A1(n2125), .A2(n2126), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .B2(n2127), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N8) );
  CLKINVX1 U2078 ( .A(n2128), .Y(n2126) );
  OAI33X1 U2079 ( .A0(n2002), .A1(n2129), .A2(n2130), .B0(n2005), .B1(n2131), 
        .B2(n2132), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N7) );
  OAI33X1 U2080 ( .A0(n2002), .A1(n2133), .A2(n2134), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .B2(n2135), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N6) );
  CLKINVX1 U2081 ( .A(n2136), .Y(n2134) );
  OAI33X1 U2082 ( .A0(n2002), .A1(n2137), .A2(n2138), .B0(n2005), .B1(n2139), 
        .B2(n2140), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N5) );
  OAI33X1 U2083 ( .A0(n2002), .A1(n2141), .A2(n2142), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .B2(n2143), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N4) );
  CLKINVX1 U2084 ( .A(n2144), .Y(n2142) );
  OAI33X1 U2085 ( .A0(n2002), .A1(n2145), .A2(n2146), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .B2(n2147), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N34) );
  CLKINVX1 U2086 ( .A(n2148), .Y(n2146) );
  OAI33X1 U2087 ( .A0(n2002), .A1(n2149), .A2(n2150), .B0(n2005), .B1(n2151), 
        .B2(n2152), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N33) );
  OAI33X1 U2088 ( .A0(n2002), .A1(n2153), .A2(n2154), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .B2(n2155), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N32) );
  CLKINVX1 U2089 ( .A(n2156), .Y(n2154) );
  OAI33X1 U2090 ( .A0(n2002), .A1(n2157), .A2(n2158), .B0(n2005), .B1(n2159), 
        .B2(n2160), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N31) );
  OAI33X1 U2091 ( .A0(n2002), .A1(n2161), .A2(n2162), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .B2(n2163), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N30) );
  CLKINVX1 U2092 ( .A(n2164), .Y(n2162) );
  OAI33X1 U2093 ( .A0(n2002), .A1(n2165), .A2(n2166), .B0(n2005), .B1(n2167), 
        .B2(n2168), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N3) );
  OAI33X1 U2094 ( .A0(n2002), .A1(n2169), .A2(n2170), .B0(n2005), .B1(n2171), 
        .B2(n2172), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N29) );
  OAI33X1 U2095 ( .A0(n2002), .A1(n2173), .A2(n2174), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .B2(n2175), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N28) );
  CLKINVX1 U2096 ( .A(n2176), .Y(n2174) );
  OAI33X1 U2097 ( .A0(n2002), .A1(n2177), .A2(n2178), .B0(n2005), .B1(n2179), 
        .B2(n2180), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N27) );
  OAI33X1 U2098 ( .A0(n2002), .A1(n2181), .A2(n2182), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .B2(n2183), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N26) );
  CLKINVX1 U2099 ( .A(n2184), .Y(n2182) );
  OAI33X1 U2100 ( .A0(n2002), .A1(n2185), .A2(n2186), .B0(n2005), .B1(n2187), 
        .B2(n2188), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N25) );
  OAI33X1 U2101 ( .A0(n2002), .A1(n2189), .A2(n2190), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .B2(n2191), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N24) );
  CLKINVX1 U2102 ( .A(n2192), .Y(n2190) );
  OAI33X1 U2103 ( .A0(n2002), .A1(n2193), .A2(n2194), .B0(n2005), .B1(n2195), 
        .B2(n2196), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N23) );
  OAI33X1 U2104 ( .A0(n2002), .A1(n2197), .A2(n2198), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .B2(n2199), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N22) );
  CLKINVX1 U2105 ( .A(n2200), .Y(n2198) );
  OAI33X1 U2106 ( .A0(n2002), .A1(n2201), .A2(n2202), .B0(n2005), .B1(n2203), 
        .B2(n2204), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N21) );
  OAI33X1 U2107 ( .A0(n2002), .A1(n2205), .A2(n2206), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .B2(n2207), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N20) );
  CLKINVX1 U2108 ( .A(n2208), .Y(n2206) );
  OAI33X1 U2109 ( .A0(n2002), .A1(n2209), .A2(n2210), .B0(n2005), .B1(n2211), 
        .B2(n2212), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N19) );
  OAI33X1 U2110 ( .A0(n2002), .A1(n2213), .A2(n2214), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .B2(n2215), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N18) );
  OAI33X1 U2111 ( .A0(n2002), .A1(n2216), .A2(n2217), .B0(n2005), .B1(n2218), 
        .B2(n2219), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N17) );
  OAI33X1 U2112 ( .A0(n2002), .A1(n2220), .A2(n2221), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .B2(n2222), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N16) );
  OAI33X1 U2113 ( .A0(n2002), .A1(n2223), .A2(n2224), .B0(n2005), .B1(n2225), 
        .B2(n2226), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N15) );
  OAI33X1 U2114 ( .A0(n2002), .A1(n2227), .A2(n2228), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .B2(n2229), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N14) );
  OAI33X1 U2115 ( .A0(n2002), .A1(n2230), .A2(n2231), .B0(n2005), .B1(n2232), 
        .B2(n2233), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N13) );
  OAI33X1 U2116 ( .A0(n2002), .A1(n2234), .A2(n2235), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .B2(n2236), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N12) );
  OAI33X1 U2117 ( .A0(n2002), .A1(n2237), .A2(n2238), .B0(n2005), .B1(n2239), 
        .B2(n2240), .Y(Inst_forkAE_CipherInst_RF_RS_EX1_N11) );
  OAI33X1 U2118 ( .A0(n2002), .A1(n2241), .A2(n2242), .B0(n2005), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .B2(n2243), .Y(
        Inst_forkAE_CipherInst_RF_RS_EX1_N10) );
  CLKINVX1 U2119 ( .A(n2245), .Y(n2242) );
  CLKNAND2X2 U2120 ( .A(n1989), .B(Inst_forkAE_CipherInst_CL_n34), .Y(n2002)
         );
  OAI221X1 U2121 ( .A0(n690), .A1(n177), .B0(n2246), .B1(n145), .C0(n2247), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_99_N3) );
  AOI22XL U2122 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_99_), 
        .B0(n236), .B1(Input2[99]), .Y(n2247) );
  CLKINVX1 U2123 ( .A(n1117), .Y(n2246) );
  CLKINVX1 U2124 ( .A(n691), .Y(n690) );
  OAI2B2X1 U2125 ( .A1N(Output2[99]), .A0(n2250), .B0(n2251), .B1(n2252), .Y(
        n691) );
  XOR2X1 U2126 ( .A(n1117), .B(n2253), .Y(Output2[99]) );
  NOR2X1 U2127 ( .A(n250), .B(n2251), .Y(n2253) );
  CLKINVX1 U2128 ( .A(Input2[99]), .Y(n2251) );
  OAI2B11X1 U2129 ( .A1N(Inst_forkAE_CipherInst_RF_S_MID_D2[98]), .A0(n2255), 
        .B0(n2256), .C0(n2257), .Y(n1117) );
  AOI22XL U2130 ( .A0(n2258), .A1(n2259), .B0(n260), .B1(n2261), .Y(n2257) );
  XOR2X1 U2131 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .B(n2262), .Y(
        n2261) );
  XOR2X1 U2132 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[66]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_18_), .Y(n2259) );
  MXI2X1 U2133 ( .A(n2263), .B(n2264), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[100]), .Y(n2256) );
  OAI21X1 U2134 ( .A0(n2265), .A1(n281), .B0(n2267), .Y(n2264) );
  NOR2X1 U2135 ( .A(n2056), .B(n2175), .Y(n2265) );
  NOR3X1 U2136 ( .A(n2175), .B(n276), .C(n2056), .Y(n2263) );
  OAI221X1 U2137 ( .A0(n694), .A1(n178), .B0(n2268), .B1(n152), .C0(n2269), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_98_N3) );
  AOI22XL U2138 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_98_), 
        .B0(n236), .B1(Input2[98]), .Y(n2269) );
  CLKINVX1 U2139 ( .A(n1119), .Y(n2268) );
  CLKINVX1 U2140 ( .A(n695), .Y(n694) );
  OAI2B2X1 U2141 ( .A1N(Output2[98]), .A0(n2250), .B0(n2270), .B1(n2252), .Y(
        n695) );
  XOR2X1 U2142 ( .A(n1119), .B(n2271), .Y(Output2[98]) );
  NOR2X1 U2143 ( .A(n245), .B(n2270), .Y(n2271) );
  CLKINVX1 U2144 ( .A(Input2[98]), .Y(n2270) );
  OAI221X1 U2145 ( .A0(n2272), .A1(n2273), .B0(n2054), .B1(n2274), .C0(n2275), 
        .Y(n1119) );
  MXI2X1 U2146 ( .A(n2276), .B(n2277), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[96]), .Y(n2275) );
  OAI21X1 U2147 ( .A0(n2278), .A1(n280), .B0(n2267), .Y(n2277) );
  NOR2X1 U2148 ( .A(n2060), .B(n2179), .Y(n2278) );
  NOR3X1 U2149 ( .A(n2266), .B(n2060), .C(n2179), .Y(n2276) );
  XOR2X1 U2150 ( .A(n2279), .B(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]), .Y(
        n2272) );
  OAI221X1 U2151 ( .A0(n698), .A1(n179), .B0(n1120), .B1(n152), .C0(n2280), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_97_N3) );
  AOI22XL U2152 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_97_), 
        .B0(n236), .B1(Input2[97]), .Y(n2280) );
  CLKINVX1 U2153 ( .A(n699), .Y(n698) );
  OAI2B2X1 U2154 ( .A1N(Output2[97]), .A0(n2250), .B0(n2281), .B1(n2252), .Y(
        n699) );
  CLKINVX1 U2155 ( .A(Input2[97]), .Y(n2281) );
  XOR2X1 U2156 ( .A(n2282), .B(n1120), .Y(Output2[97]) );
  CLKINVX1 U2157 ( .A(n2283), .Y(n1120) );
  OAI221X1 U2158 ( .A0(n2284), .A1(n2273), .B0(n2173), .B1(n2274), .C0(n2285), 
        .Y(n2283) );
  AOI2BB2X1 U2159 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[99]), .B1(n294), 
        .A0N(n285), .A1N(n2179), .Y(n2285) );
  XOR2X1 U2160 ( .A(n2287), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[31]), .Y(
        n2284) );
  CLKNAND2X2 U2161 ( .A(Input2[97]), .B(n2288), .Y(n2282) );
  OAI221X1 U2162 ( .A0(n702), .A1(n171), .B0(n1121), .B1(n152), .C0(n2289), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_96_N3) );
  AOI22XL U2163 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_96_), 
        .B0(n235), .B1(Input2[96]), .Y(n2289) );
  CLKINVX1 U2164 ( .A(n703), .Y(n702) );
  OAI2B2X1 U2165 ( .A1N(Output2[96]), .A0(n2250), .B0(n2290), .B1(n2252), .Y(
        n703) );
  XNOR2X1 U2166 ( .A(n1121), .B(n2291), .Y(Output2[96]) );
  NOR2X1 U2167 ( .A(n245), .B(n2290), .Y(n2291) );
  CLKINVX1 U2168 ( .A(Input2[96]), .Y(n2290) );
  AOI221XL U2169 ( .A0(n2292), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C2[96]), .C0(n2294), .Y(n1121) );
  AO22X1 U2170 ( .A0(n266), .A1(n2295), .B0(n301), .B1(n2296), .Y(n2294) );
  XOR2X1 U2171 ( .A(n2297), .B(n2298), .Y(n2295) );
  CLKINVX1 U2172 ( .A(n2058), .Y(n2292) );
  OAI221X1 U2173 ( .A0(n2299), .A1(n2300), .B0(n2301), .B1(n2302), .C0(n2303), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_95_N3) );
  AOI2BB2X1 U2174 ( .B0(n183), .B1(n706), .A0N(n159), .A1N(n1122), .Y(n2303)
         );
  OAI2B2X1 U2175 ( .A1N(Output2[95]), .A0(n2304), .B0(n2301), .B1(n2305), .Y(
        n706) );
  XNOR2X1 U2176 ( .A(n1122), .B(n2306), .Y(Output2[95]) );
  NOR2X1 U2177 ( .A(n245), .B(n2301), .Y(n2306) );
  AOI221XL U2178 ( .A0(n2307), .A1(n264), .B0(n295), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .C0(n2308), .Y(n1122) );
  CLKINVX1 U2179 ( .A(n2309), .Y(n2308) );
  AOI222XL U2180 ( .A0(n287), .A1(n2310), .B0(n2258), .B1(n2311), .C0(n2312), 
        .C1(n2313), .Y(n2309) );
  XOR2X1 U2181 ( .A(n2314), .B(n2315), .Y(n2311) );
  XOR2X1 U2182 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[39]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_45_), .Y(n2315) );
  CLKINVX1 U2183 ( .A(Input2[95]), .Y(n2301) );
  CLKINVX1 U2184 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_95_), .Y(n2299) );
  OAI221X1 U2185 ( .A0(n709), .A1(n172), .B0(n1124), .B1(n152), .C0(n2316), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_94_N3) );
  AOI22XL U2186 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_94_), 
        .B0(n235), .B1(Input2[94]), .Y(n2316) );
  CLKINVX1 U2187 ( .A(n710), .Y(n709) );
  OAI2B2X1 U2188 ( .A1N(Input2[94]), .A0(n2305), .B0(n2317), .B1(n2304), .Y(
        n710) );
  CLKINVX1 U2189 ( .A(Output2[94]), .Y(n2317) );
  XOR2X1 U2190 ( .A(n2318), .B(n1124), .Y(Output2[94]) );
  AOI221XL U2191 ( .A0(n2319), .A1(n2293), .B0(n2320), .B1(n265), .C0(n2321), 
        .Y(n1124) );
  AO22X1 U2192 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[90]), .A1(n301), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .B1(n292), .Y(n2321) );
  XNOR2X1 U2193 ( .A(n2322), .B(n2323), .Y(n2319) );
  MXI2X1 U2194 ( .A(n2324), .B(n2325), .S0(n313), .Y(n2323) );
  XOR2X1 U2195 ( .A(n2326), .B(n2327), .Y(n2325) );
  XOR2X1 U2196 ( .A(n2328), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .Y(
        n2326) );
  CLKINVX1 U2197 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[92]), .Y(n2324) );
  OR2X1 U2198 ( .A(n2181), .B(n2062), .Y(n2322) );
  CLKNAND2X2 U2199 ( .A(Input2[94]), .B(n2288), .Y(n2318) );
  OAI221X1 U2200 ( .A0(n713), .A1(n173), .B0(n1125), .B1(n152), .C0(n2329), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_93_N3) );
  AOI22XL U2201 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_93_), 
        .B0(n235), .B1(Input2[93]), .Y(n2329) );
  CLKINVX1 U2202 ( .A(n714), .Y(n713) );
  OAI2B2X1 U2203 ( .A1N(Output2[93]), .A0(n2304), .B0(n2330), .B1(n2305), .Y(
        n714) );
  XNOR2X1 U2204 ( .A(n1125), .B(n2331), .Y(Output2[93]) );
  NOR2X1 U2205 ( .A(n245), .B(n2330), .Y(n2331) );
  CLKINVX1 U2206 ( .A(Input2[93]), .Y(n2330) );
  AOI222XL U2207 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D2[95]), 
        .B0(n2333), .B1(n2293), .C0(n2334), .C1(n265), .Y(n1125) );
  XNOR2X1 U2208 ( .A(n2335), .B(n2336), .Y(n2333) );
  MXI2X1 U2209 ( .A(n2337), .B(n2338), .S0(n306), .Y(n2336) );
  XOR2X1 U2210 ( .A(n2339), .B(n2340), .Y(n2338) );
  XOR2X1 U2211 ( .A(n2341), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .Y(
        n2339) );
  CLKNAND2X2 U2212 ( .A(n2342), .B(n2343), .Y(n2335) );
  OAI221X1 U2213 ( .A0(n717), .A1(n176), .B0(n1127), .B1(n152), .C0(n2344), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_92_N3) );
  AOI22XL U2214 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_92_), 
        .B0(n235), .B1(Input2[92]), .Y(n2344) );
  CLKINVX1 U2215 ( .A(n718), .Y(n717) );
  OAI2B2X1 U2216 ( .A1N(Input2[92]), .A0(n2305), .B0(n2345), .B1(n2304), .Y(
        n718) );
  CLKINVX1 U2217 ( .A(Output2[92]), .Y(n2345) );
  XOR2X1 U2218 ( .A(n2346), .B(n1127), .Y(Output2[92]) );
  AOI221XL U2219 ( .A0(n2347), .A1(n295), .B0(n2343), .B1(n2293), .C0(n2348), 
        .Y(n1127) );
  OAI2BB2X1 U2220 ( .B0(n2064), .B1(n285), .A0N(n2349), .A1N(n269), .Y(n2348)
         );
  CLKINVX1 U2221 ( .A(n2185), .Y(n2343) );
  MXI2X1 U2222 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[91]), .B(n2350), .S0(
        n306), .Y(n2185) );
  XOR2X1 U2223 ( .A(n2351), .B(n2352), .Y(n2350) );
  XOR2X1 U2224 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[51]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_43_), .Y(n2352) );
  CLKNAND2X2 U2225 ( .A(Input2[92]), .B(n2288), .Y(n2346) );
  OAI221X1 U2226 ( .A0(n721), .A1(n174), .B0(n2353), .B1(n152), .C0(n2354), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_91_N3) );
  AOI22XL U2227 ( .A0(n208), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_91_), 
        .B0(n235), .B1(Input2[91]), .Y(n2354) );
  CLKINVX1 U2228 ( .A(n1129), .Y(n2353) );
  CLKINVX1 U2229 ( .A(n722), .Y(n721) );
  OAI2B2X1 U2230 ( .A1N(Output2[91]), .A0(n2304), .B0(n2355), .B1(n2305), .Y(
        n722) );
  XOR2X1 U2231 ( .A(n1129), .B(n2356), .Y(Output2[91]) );
  NOR2X1 U2232 ( .A(n245), .B(n2355), .Y(n2356) );
  CLKINVX1 U2233 ( .A(Input2[91]), .Y(n2355) );
  OAI2B11X1 U2234 ( .A1N(n2357), .A0(n2273), .B0(n2358), .C0(n2359), .Y(n1129)
         );
  AOI22XL U2235 ( .A0(n2258), .A1(n2360), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[90]), .B1(n2312), .Y(n2359) );
  XNOR2X1 U2236 ( .A(n2361), .B(n2362), .Y(n2360) );
  XOR2X1 U2237 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[50]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_42_), .Y(n2362) );
  MXI2X1 U2238 ( .A(n2363), .B(n2364), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[92]), .Y(n2358) );
  OAI21X1 U2239 ( .A0(n2365), .A1(n280), .B0(n2267), .Y(n2364) );
  NOR2X1 U2240 ( .A(n2064), .B(n2183), .Y(n2365) );
  NOR3X1 U2241 ( .A(n2183), .B(n276), .C(n2064), .Y(n2363) );
  CLKINVX1 U2242 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[92]), .Y(n2064) );
  CLKINVX1 U2243 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[95]), .Y(n2183) );
  OAI221X1 U2244 ( .A0(n725), .A1(n172), .B0(n1130), .B1(n152), .C0(n2366), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_90_N3) );
  AOI22XL U2245 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_90_), 
        .B0(n235), .B1(Input2[90]), .Y(n2366) );
  CLKINVX1 U2246 ( .A(n726), .Y(n725) );
  OAI2B2X1 U2247 ( .A1N(Output2[90]), .A0(n2304), .B0(n2367), .B1(n2305), .Y(
        n726) );
  XNOR2X1 U2248 ( .A(n1130), .B(n2368), .Y(Output2[90]) );
  NOR2X1 U2249 ( .A(n245), .B(n2367), .Y(n2368) );
  CLKINVX1 U2250 ( .A(Input2[90]), .Y(n2367) );
  AOI221XL U2251 ( .A0(n2369), .A1(n2293), .B0(n2370), .B1(n265), .C0(n2371), 
        .Y(n1130) );
  MX2X1 U2252 ( .A(n2372), .B(n2373), .S0(n2337), .Y(n2371) );
  CLKINVX1 U2253 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[88]), .Y(n2337) );
  NOR3X1 U2254 ( .A(n2266), .B(n2067), .C(n2187), .Y(n2373) );
  OAI21X1 U2255 ( .A0(n2374), .A1(n279), .B0(n2267), .Y(n2372) );
  NOR2X1 U2256 ( .A(n2067), .B(n2187), .Y(n2374) );
  CLKINVX1 U2257 ( .A(n2062), .Y(n2369) );
  MXI2X1 U2258 ( .A(n2347), .B(n2375), .S0(n306), .Y(n2062) );
  XOR2X1 U2259 ( .A(n2376), .B(n2377), .Y(n2375) );
  XOR2X1 U2260 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[34]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_), .Y(n2377) );
  XOR2X1 U2261 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_23_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[92]), .Y(n2347) );
  OAI221X1 U2262 ( .A0(n1039), .A1(n173), .B0(n1268), .B1(n152), .C0(n2378), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_9_N3) );
  AOI22XL U2263 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_9_), 
        .B0(n235), .B1(Input2[9]), .Y(n2378) );
  CLKINVX1 U2264 ( .A(n1040), .Y(n1039) );
  OAI2B2X1 U2265 ( .A1N(Output2[9]), .A0(n2379), .B0(n2380), .B1(n2381), .Y(
        n1040) );
  CLKINVX1 U2266 ( .A(Input2[9]), .Y(n2380) );
  XOR2X1 U2267 ( .A(n2382), .B(n1268), .Y(Output2[9]) );
  CLKINVX1 U2268 ( .A(n2383), .Y(n1268) );
  OAI221X1 U2269 ( .A0(n2133), .A1(n2274), .B0(n2384), .B1(n2273), .C0(n2385), 
        .Y(n2383) );
  AOI22XL U2270 ( .A0(n291), .A1(n2386), .B0(n294), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D2[11]), .Y(n2385) );
  CLKNAND2X2 U2271 ( .A(Input2[9]), .B(n2288), .Y(n2382) );
  OAI221X1 U2272 ( .A0(n729), .A1(n176), .B0(n2387), .B1(n152), .C0(n2388), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_89_N3) );
  AOI22XL U2273 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_89_), 
        .B0(n235), .B1(Input2[89]), .Y(n2388) );
  CLKINVX1 U2274 ( .A(n1132), .Y(n2387) );
  CLKINVX1 U2275 ( .A(n730), .Y(n729) );
  OAI2B2X1 U2276 ( .A1N(Output2[89]), .A0(n2304), .B0(n2389), .B1(n2305), .Y(
        n730) );
  XOR2X1 U2277 ( .A(n1132), .B(n2390), .Y(Output2[89]) );
  NOR2X1 U2278 ( .A(n245), .B(n2389), .Y(n2390) );
  CLKINVX1 U2279 ( .A(Input2[89]), .Y(n2389) );
  OAI221X1 U2280 ( .A0(n2181), .A1(n2274), .B0(n2187), .B1(n278), .C0(n2391), 
        .Y(n1132) );
  AOI22XL U2281 ( .A0(n261), .A1(n2392), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[91]), .B1(n300), .Y(n2391) );
  MXI2X1 U2282 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[95]), .B(n2393), .S0(
        n306), .Y(n2181) );
  XOR2X1 U2283 ( .A(n2394), .B(n2395), .Y(n2393) );
  XOR2X1 U2284 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[55]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_47_), .Y(n2395) );
  OAI221X1 U2285 ( .A0(n733), .A1(n174), .B0(n1134), .B1(n152), .C0(n2396), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_88_N3) );
  AOI22XL U2286 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_88_), 
        .B0(n235), .B1(Input2[88]), .Y(n2396) );
  CLKINVX1 U2287 ( .A(n734), .Y(n733) );
  OAI2B2X1 U2288 ( .A1N(Input2[88]), .A0(n2305), .B0(n2397), .B1(n2304), .Y(
        n734) );
  CLKINVX1 U2289 ( .A(Output2[88]), .Y(n2397) );
  XOR2X1 U2290 ( .A(n2398), .B(n1134), .Y(Output2[88]) );
  AOI221XL U2291 ( .A0(n2313), .A1(n296), .B0(n2342), .B1(n2293), .C0(n2399), 
        .Y(n1134) );
  AO22X1 U2292 ( .A0(n266), .A1(n2400), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C2[88]), .B1(n292), .Y(n2399) );
  CLKINVX1 U2293 ( .A(n2065), .Y(n2342) );
  MXI2X1 U2294 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .B(n2401), .S0(
        n306), .Y(n2065) );
  XOR2X1 U2295 ( .A(n2402), .B(n2403), .Y(n2401) );
  XOR2X1 U2296 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[49]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_41_), .Y(n2403) );
  XOR2X1 U2297 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_22_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[88]), .Y(n2313) );
  CLKNAND2X2 U2298 ( .A(Input2[88]), .B(n2288), .Y(n2398) );
  OAI221X1 U2299 ( .A0(n2404), .A1(n2300), .B0(n2405), .B1(n2302), .C0(n2406), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_87_N3) );
  AOI2BB2X1 U2300 ( .B0(n181), .B1(n737), .A0N(n159), .A1N(n1135), .Y(n2406)
         );
  OAI2B2X1 U2301 ( .A1N(Output2[87]), .A0(n2407), .B0(n2405), .B1(n2408), .Y(
        n737) );
  XNOR2X1 U2302 ( .A(n1135), .B(n2409), .Y(Output2[87]) );
  NOR2X1 U2303 ( .A(n245), .B(n2405), .Y(n2409) );
  AOI221XL U2304 ( .A0(n2410), .A1(n264), .B0(n295), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .C0(n2411), .Y(n1135) );
  CLKINVX1 U2305 ( .A(n2412), .Y(n2411) );
  AOI222XL U2306 ( .A0(n288), .A1(n2413), .B0(n2258), .B1(n2414), .C0(n2312), 
        .C1(n2415), .Y(n2412) );
  XOR2X1 U2307 ( .A(n2416), .B(n2417), .Y(n2414) );
  XOR2X1 U2308 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[63]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_13_), .Y(n2417) );
  CLKINVX1 U2309 ( .A(Input2[87]), .Y(n2405) );
  CLKINVX1 U2310 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_87_), .Y(n2404) );
  OAI221X1 U2311 ( .A0(n740), .A1(n175), .B0(n1137), .B1(n151), .C0(n2418), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_86_N3) );
  AOI22XL U2312 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_86_), 
        .B0(n235), .B1(Input2[86]), .Y(n2418) );
  CLKINVX1 U2313 ( .A(n741), .Y(n740) );
  OAI2B2X1 U2314 ( .A1N(Input2[86]), .A0(n2408), .B0(n2419), .B1(n2407), .Y(
        n741) );
  CLKINVX1 U2315 ( .A(Output2[86]), .Y(n2419) );
  XOR2X1 U2316 ( .A(n2420), .B(n1137), .Y(Output2[86]) );
  AOI221XL U2317 ( .A0(n2421), .A1(n2293), .B0(n2422), .B1(n265), .C0(n2423), 
        .Y(n1137) );
  AO22X1 U2318 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[82]), .A1(n301), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .B1(n292), .Y(n2423) );
  XNOR2X1 U2319 ( .A(n2424), .B(n2425), .Y(n2421) );
  MXI2X1 U2320 ( .A(n2426), .B(n2427), .S0(n306), .Y(n2425) );
  XOR2X1 U2321 ( .A(n2428), .B(n2429), .Y(n2427) );
  XOR2X1 U2322 ( .A(n2430), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[44]), .Y(
        n2428) );
  CLKINVX1 U2323 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[84]), .Y(n2426) );
  OR2X1 U2324 ( .A(n2189), .B(n2069), .Y(n2424) );
  CLKNAND2X2 U2325 ( .A(Input2[86]), .B(n2288), .Y(n2420) );
  OAI221X1 U2326 ( .A0(n744), .A1(n168), .B0(n1138), .B1(n151), .C0(n2431), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_85_N3) );
  AOI22XL U2327 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_85_), 
        .B0(n235), .B1(Input2[85]), .Y(n2431) );
  CLKINVX1 U2328 ( .A(n745), .Y(n744) );
  OAI2B2X1 U2329 ( .A1N(Output2[85]), .A0(n2407), .B0(n2432), .B1(n2408), .Y(
        n745) );
  XNOR2X1 U2330 ( .A(n1138), .B(n2433), .Y(Output2[85]) );
  NOR2X1 U2331 ( .A(n245), .B(n2432), .Y(n2433) );
  CLKINVX1 U2332 ( .A(Input2[85]), .Y(n2432) );
  AOI222XL U2333 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D2[87]), 
        .B0(n2434), .B1(n2293), .C0(n2435), .C1(n265), .Y(n1138) );
  XNOR2X1 U2334 ( .A(n2436), .B(n2437), .Y(n2434) );
  MXI2X1 U2335 ( .A(n2438), .B(n2439), .S0(n306), .Y(n2437) );
  XOR2X1 U2336 ( .A(n2440), .B(n2441), .Y(n2439) );
  XOR2X1 U2337 ( .A(n2442), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[40]), .Y(
        n2440) );
  CLKNAND2X2 U2338 ( .A(n2443), .B(n2444), .Y(n2436) );
  OAI221X1 U2339 ( .A0(n748), .A1(n169), .B0(n1140), .B1(n151), .C0(n2445), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_84_N3) );
  AOI22XL U2340 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_84_), 
        .B0(n235), .B1(Input2[84]), .Y(n2445) );
  CLKINVX1 U2341 ( .A(n749), .Y(n748) );
  OAI2B2X1 U2342 ( .A1N(Input2[84]), .A0(n2408), .B0(n2446), .B1(n2407), .Y(
        n749) );
  CLKINVX1 U2343 ( .A(Output2[84]), .Y(n2446) );
  XOR2X1 U2344 ( .A(n2447), .B(n1140), .Y(Output2[84]) );
  AOI221XL U2345 ( .A0(n2448), .A1(n296), .B0(n2444), .B1(n2293), .C0(n2449), 
        .Y(n1140) );
  OAI2BB2X1 U2346 ( .B0(n2071), .B1(n284), .A0N(n2450), .A1N(n269), .Y(n2449)
         );
  CLKINVX1 U2347 ( .A(n2193), .Y(n2444) );
  MXI2X1 U2348 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[83]), .B(n2451), .S0(
        n306), .Y(n2193) );
  XOR2X1 U2349 ( .A(n2452), .B(n2453), .Y(n2451) );
  XOR2X1 U2350 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[43]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_11_), .Y(n2453) );
  CLKNAND2X2 U2351 ( .A(Input2[84]), .B(n2288), .Y(n2447) );
  OAI221X1 U2352 ( .A0(n752), .A1(n170), .B0(n2454), .B1(n151), .C0(n2455), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_83_N3) );
  AOI22XL U2353 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_83_), 
        .B0(n235), .B1(Input2[83]), .Y(n2455) );
  CLKINVX1 U2354 ( .A(n1142), .Y(n2454) );
  CLKINVX1 U2355 ( .A(n753), .Y(n752) );
  OAI2B2X1 U2356 ( .A1N(Output2[83]), .A0(n2407), .B0(n2456), .B1(n2408), .Y(
        n753) );
  XOR2X1 U2357 ( .A(n1142), .B(n2457), .Y(Output2[83]) );
  NOR2X1 U2358 ( .A(n245), .B(n2456), .Y(n2457) );
  CLKINVX1 U2359 ( .A(Input2[83]), .Y(n2456) );
  OAI2B11X1 U2360 ( .A1N(n2458), .A0(n2273), .B0(n2459), .C0(n2460), .Y(n1142)
         );
  AOI22XL U2361 ( .A0(n2258), .A1(n2461), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[82]), .B1(n2312), .Y(n2460) );
  XNOR2X1 U2362 ( .A(n2462), .B(n2463), .Y(n2461) );
  XOR2X1 U2363 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[42]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_10_), .Y(n2463) );
  MXI2X1 U2364 ( .A(n2464), .B(n2465), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[84]), .Y(n2459) );
  OAI21X1 U2365 ( .A0(n2466), .A1(n280), .B0(n2267), .Y(n2465) );
  NOR2X1 U2366 ( .A(n2071), .B(n2191), .Y(n2466) );
  NOR3X1 U2367 ( .A(n2191), .B(n276), .C(n2071), .Y(n2464) );
  CLKINVX1 U2368 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[84]), .Y(n2071) );
  CLKINVX1 U2369 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[87]), .Y(n2191) );
  OAI221X1 U2370 ( .A0(n756), .A1(n167), .B0(n1143), .B1(n151), .C0(n2467), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_82_N3) );
  AOI22XL U2371 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_82_), 
        .B0(n234), .B1(Input2[82]), .Y(n2467) );
  CLKINVX1 U2372 ( .A(n757), .Y(n756) );
  OAI2B2X1 U2373 ( .A1N(Output2[82]), .A0(n2407), .B0(n2468), .B1(n2408), .Y(
        n757) );
  XNOR2X1 U2374 ( .A(n1143), .B(n2469), .Y(Output2[82]) );
  NOR2X1 U2375 ( .A(n245), .B(n2468), .Y(n2469) );
  CLKINVX1 U2376 ( .A(Input2[82]), .Y(n2468) );
  AOI221XL U2377 ( .A0(n2470), .A1(n2293), .B0(n2471), .B1(n266), .C0(n2472), 
        .Y(n1143) );
  MX2X1 U2378 ( .A(n2473), .B(n2474), .S0(n2438), .Y(n2472) );
  CLKINVX1 U2379 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[80]), .Y(n2438) );
  NOR3X1 U2380 ( .A(n2266), .B(n2074), .C(n2195), .Y(n2474) );
  OAI21X1 U2381 ( .A0(n2475), .A1(n279), .B0(n2267), .Y(n2473) );
  NOR2X1 U2382 ( .A(n2074), .B(n2195), .Y(n2475) );
  CLKINVX1 U2383 ( .A(n2069), .Y(n2470) );
  MXI2X1 U2384 ( .A(n2448), .B(n2476), .S0(n306), .Y(n2069) );
  XOR2X1 U2385 ( .A(n2477), .B(n2478), .Y(n2476) );
  XOR2X1 U2386 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[58]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_14_), .Y(n2478) );
  XOR2X1 U2387 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_21_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[84]), .Y(n2448) );
  OAI221X1 U2388 ( .A0(n760), .A1(n177), .B0(n2479), .B1(n151), .C0(n2480), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_81_N3) );
  AOI22XL U2389 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_81_), 
        .B0(n234), .B1(Input2[81]), .Y(n2480) );
  CLKINVX1 U2390 ( .A(n1145), .Y(n2479) );
  CLKINVX1 U2391 ( .A(n761), .Y(n760) );
  OAI2B2X1 U2392 ( .A1N(Output2[81]), .A0(n2407), .B0(n2481), .B1(n2408), .Y(
        n761) );
  XOR2X1 U2393 ( .A(n1145), .B(n2482), .Y(Output2[81]) );
  NOR2X1 U2394 ( .A(n245), .B(n2481), .Y(n2482) );
  CLKINVX1 U2395 ( .A(Input2[81]), .Y(n2481) );
  OAI221X1 U2396 ( .A0(n2189), .A1(n2274), .B0(n2195), .B1(n278), .C0(n2483), 
        .Y(n1145) );
  AOI22XL U2397 ( .A0(n261), .A1(n2484), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[83]), .B1(n300), .Y(n2483) );
  MXI2X1 U2398 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[87]), .B(n2485), .S0(
        n306), .Y(n2189) );
  XOR2X1 U2399 ( .A(n2486), .B(n2487), .Y(n2485) );
  XOR2X1 U2400 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[47]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_15_), .Y(n2487) );
  OAI221X1 U2401 ( .A0(n764), .A1(n166), .B0(n1147), .B1(n151), .C0(n2488), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_80_N3) );
  AOI22XL U2402 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_80_), 
        .B0(n234), .B1(Input2[80]), .Y(n2488) );
  CLKINVX1 U2403 ( .A(n765), .Y(n764) );
  OAI2B2X1 U2404 ( .A1N(Input2[80]), .A0(n2408), .B0(n2489), .B1(n2407), .Y(
        n765) );
  CLKINVX1 U2405 ( .A(Output2[80]), .Y(n2489) );
  XOR2X1 U2406 ( .A(n2490), .B(n1147), .Y(Output2[80]) );
  AOI221XL U2407 ( .A0(n2415), .A1(n296), .B0(n2443), .B1(n2293), .C0(n2491), 
        .Y(n1147) );
  AO22X1 U2408 ( .A0(n266), .A1(n2492), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C2[80]), .B1(n292), .Y(n2491) );
  CLKINVX1 U2409 ( .A(n2072), .Y(n2443) );
  MXI2X1 U2410 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .B(n2493), .S0(
        n306), .Y(n2072) );
  XOR2X1 U2411 ( .A(n2494), .B(n2495), .Y(n2493) );
  XOR2X1 U2412 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[41]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_9_), .Y(n2495) );
  XOR2X1 U2413 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_20_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[80]), .Y(n2415) );
  CLKNAND2X2 U2414 ( .A(Input2[80]), .B(n2288), .Y(n2490) );
  OAI221X1 U2415 ( .A0(n1043), .A1(n165), .B0(n1270), .B1(n151), .C0(n2496), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_8_N3) );
  AOI22XL U2416 ( .A0(n207), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_8_), 
        .B0(n234), .B1(Input2[8]), .Y(n2496) );
  CLKINVX1 U2417 ( .A(n1044), .Y(n1043) );
  OAI2B2X1 U2418 ( .A1N(Input2[8]), .A0(n2381), .B0(n2497), .B1(n2379), .Y(
        n1044) );
  CLKINVX1 U2419 ( .A(Output2[8]), .Y(n2497) );
  XOR2X1 U2420 ( .A(n2498), .B(n1270), .Y(Output2[8]) );
  AOI221XL U2421 ( .A0(n2499), .A1(n296), .B0(n2500), .B1(n2293), .C0(n2501), 
        .Y(n1270) );
  OAI2BB2X1 U2422 ( .B0(n2502), .B1(n284), .A0N(n2503), .A1N(n269), .Y(n2501)
         );
  CLKNAND2X2 U2423 ( .A(Input2[8]), .B(n2288), .Y(n2498) );
  OAI221X1 U2424 ( .A0(n2504), .A1(n2300), .B0(n2505), .B1(n2302), .C0(n2506), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_79_N3) );
  AOI22XL U2425 ( .A0(n185), .A1(n768), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1149), .Y(n2506) );
  OAI2B2X1 U2426 ( .A1N(Output2[79]), .A0(n2507), .B0(n2505), .B1(n2508), .Y(
        n768) );
  XOR2X1 U2427 ( .A(n1149), .B(n2509), .Y(Output2[79]) );
  NOR2X1 U2428 ( .A(n245), .B(n2505), .Y(n2509) );
  OAI221X1 U2429 ( .A0(n2510), .A1(n2273), .B0(n2267), .B1(n2511), .C0(n2512), 
        .Y(n1149) );
  AOI222XL U2430 ( .A0(n289), .A1(n2513), .B0(n2258), .B1(n2514), .C0(n2312), 
        .C1(n2515), .Y(n2512) );
  XOR2X1 U2431 ( .A(n2516), .B(n2517), .Y(n2514) );
  XOR2X1 U2432 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[55]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_29_), .Y(n2517) );
  CLKINVX1 U2433 ( .A(n2518), .Y(n2510) );
  CLKINVX1 U2434 ( .A(Input2[79]), .Y(n2505) );
  CLKINVX1 U2435 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_79_), .Y(n2504) );
  OAI221X1 U2436 ( .A0(n771), .A1(n175), .B0(n1151), .B1(n151), .C0(n2519), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_78_N3) );
  AOI22XL U2437 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_78_), 
        .B0(n234), .B1(Input2[78]), .Y(n2519) );
  CLKINVX1 U2438 ( .A(n772), .Y(n771) );
  OAI2B2X1 U2439 ( .A1N(Input2[78]), .A0(n2508), .B0(n2520), .B1(n2507), .Y(
        n772) );
  CLKINVX1 U2440 ( .A(Output2[78]), .Y(n2520) );
  XOR2X1 U2441 ( .A(n2521), .B(n1151), .Y(Output2[78]) );
  AOI221XL U2442 ( .A0(n2522), .A1(n2293), .B0(n2523), .B1(n265), .C0(n2524), 
        .Y(n1151) );
  OAI2BB2X1 U2443 ( .B0(n2511), .B1(n284), .A0N(
        Inst_forkAE_CipherInst_RF_S_MID_D2[74]), .A1N(n301), .Y(n2524) );
  CLKINVX1 U2444 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[73]), .Y(n2511) );
  XNOR2X1 U2445 ( .A(n2525), .B(n2526), .Y(n2522) );
  MXI2X1 U2446 ( .A(n2527), .B(n2528), .S0(n307), .Y(n2526) );
  XOR2X1 U2447 ( .A(n2529), .B(n2530), .Y(n2528) );
  XOR2X1 U2448 ( .A(n2531), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[36]), .Y(
        n2529) );
  CLKINVX1 U2449 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[76]), .Y(n2527) );
  OR2X1 U2450 ( .A(n2197), .B(n2076), .Y(n2525) );
  CLKNAND2X2 U2451 ( .A(Input2[78]), .B(n2288), .Y(n2521) );
  OAI221X1 U2452 ( .A0(n775), .A1(n168), .B0(n1152), .B1(n151), .C0(n2532), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_77_N3) );
  AOI22XL U2453 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_77_), 
        .B0(n234), .B1(Input2[77]), .Y(n2532) );
  CLKINVX1 U2454 ( .A(n776), .Y(n775) );
  OAI2B2X1 U2455 ( .A1N(Output2[77]), .A0(n2507), .B0(n2533), .B1(n2508), .Y(
        n776) );
  XNOR2X1 U2456 ( .A(n1152), .B(n2534), .Y(Output2[77]) );
  NOR2X1 U2457 ( .A(n245), .B(n2533), .Y(n2534) );
  CLKINVX1 U2458 ( .A(Input2[77]), .Y(n2533) );
  AOI222XL U2459 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D2[79]), 
        .B0(n2535), .B1(n2293), .C0(n2536), .C1(n265), .Y(n1152) );
  XNOR2X1 U2460 ( .A(n2537), .B(n2538), .Y(n2535) );
  MXI2X1 U2461 ( .A(n2539), .B(n2540), .S0(n307), .Y(n2538) );
  XOR2X1 U2462 ( .A(n2541), .B(n2542), .Y(n2540) );
  XOR2X1 U2463 ( .A(n2543), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[32]), .Y(
        n2541) );
  CLKNAND2X2 U2464 ( .A(n2544), .B(n2545), .Y(n2537) );
  OAI221X1 U2465 ( .A0(n779), .A1(n169), .B0(n1154), .B1(n151), .C0(n2546), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_76_N3) );
  AOI22XL U2466 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_76_), 
        .B0(n234), .B1(Input2[76]), .Y(n2546) );
  CLKINVX1 U2467 ( .A(n780), .Y(n779) );
  OAI2B2X1 U2468 ( .A1N(Input2[76]), .A0(n2508), .B0(n2547), .B1(n2507), .Y(
        n780) );
  CLKINVX1 U2469 ( .A(Output2[76]), .Y(n2547) );
  XOR2X1 U2470 ( .A(n2548), .B(n1154), .Y(Output2[76]) );
  AOI221XL U2471 ( .A0(n2549), .A1(n296), .B0(n2545), .B1(n2293), .C0(n2550), 
        .Y(n1154) );
  OAI2BB2X1 U2472 ( .B0(n2078), .B1(n284), .A0N(n2551), .A1N(n268), .Y(n2550)
         );
  CLKINVX1 U2473 ( .A(n2201), .Y(n2545) );
  MXI2X1 U2474 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[75]), .B(n2552), .S0(
        n307), .Y(n2201) );
  XOR2X1 U2475 ( .A(n2553), .B(n2554), .Y(n2552) );
  XOR2X1 U2476 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[35]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_27_), .Y(n2554) );
  CLKNAND2X2 U2477 ( .A(Input2[76]), .B(n2288), .Y(n2548) );
  OAI221X1 U2478 ( .A0(n783), .A1(n170), .B0(n2555), .B1(n151), .C0(n2556), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_75_N3) );
  AOI22XL U2479 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_75_), 
        .B0(n234), .B1(Input2[75]), .Y(n2556) );
  CLKINVX1 U2480 ( .A(n1156), .Y(n2555) );
  CLKINVX1 U2481 ( .A(n784), .Y(n783) );
  OAI2B2X1 U2482 ( .A1N(Output2[75]), .A0(n2507), .B0(n2557), .B1(n2508), .Y(
        n784) );
  XOR2X1 U2483 ( .A(n1156), .B(n2558), .Y(Output2[75]) );
  NOR2X1 U2484 ( .A(n246), .B(n2557), .Y(n2558) );
  CLKINVX1 U2485 ( .A(Input2[75]), .Y(n2557) );
  OAI2B11X1 U2486 ( .A1N(n2559), .A0(n2273), .B0(n2560), .C0(n2561), .Y(n1156)
         );
  AOI22XL U2487 ( .A0(n2258), .A1(n2562), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[74]), .B1(n2312), .Y(n2561) );
  XNOR2X1 U2488 ( .A(n2563), .B(n2564), .Y(n2562) );
  XOR2X1 U2489 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[34]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_26_), .Y(n2564) );
  MXI2X1 U2490 ( .A(n2565), .B(n2566), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[76]), .Y(n2560) );
  OAI21X1 U2491 ( .A0(n2567), .A1(n279), .B0(n2267), .Y(n2566) );
  NOR2X1 U2492 ( .A(n2078), .B(n2199), .Y(n2567) );
  NOR3X1 U2493 ( .A(n2199), .B(n276), .C(n2078), .Y(n2565) );
  CLKINVX1 U2494 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[76]), .Y(n2078) );
  CLKINVX1 U2495 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[79]), .Y(n2199) );
  OAI221X1 U2496 ( .A0(n787), .A1(n167), .B0(n1157), .B1(n151), .C0(n2568), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_74_N3) );
  AOI22XL U2497 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_74_), 
        .B0(n234), .B1(Input2[74]), .Y(n2568) );
  CLKINVX1 U2498 ( .A(n788), .Y(n787) );
  OAI2B2X1 U2499 ( .A1N(Output2[74]), .A0(n2507), .B0(n2569), .B1(n2508), .Y(
        n788) );
  XNOR2X1 U2500 ( .A(n1157), .B(n2570), .Y(Output2[74]) );
  NOR2X1 U2501 ( .A(n246), .B(n2569), .Y(n2570) );
  CLKINVX1 U2502 ( .A(Input2[74]), .Y(n2569) );
  AOI221XL U2503 ( .A0(n2571), .A1(n2293), .B0(n2572), .B1(n266), .C0(n2573), 
        .Y(n1157) );
  MX2X1 U2504 ( .A(n2574), .B(n2575), .S0(n2539), .Y(n2573) );
  NOR3X1 U2505 ( .A(n280), .B(n2081), .C(n2203), .Y(n2575) );
  OAI21X1 U2506 ( .A0(n2576), .A1(n279), .B0(n2267), .Y(n2574) );
  NOR2X1 U2507 ( .A(n2081), .B(n2203), .Y(n2576) );
  CLKINVX1 U2508 ( .A(n2076), .Y(n2571) );
  MXI2X1 U2509 ( .A(n2549), .B(n2577), .S0(n307), .Y(n2076) );
  XOR2X1 U2510 ( .A(n2578), .B(n2579), .Y(n2577) );
  XOR2X1 U2511 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[50]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_), .Y(n2579) );
  XOR2X1 U2512 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_19_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[76]), .Y(n2549) );
  OAI221X1 U2513 ( .A0(n791), .A1(n178), .B0(n2580), .B1(n151), .C0(n2581), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_73_N3) );
  AOI22XL U2514 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_73_), 
        .B0(n234), .B1(Input2[73]), .Y(n2581) );
  CLKINVX1 U2515 ( .A(n1159), .Y(n2580) );
  CLKINVX1 U2516 ( .A(n792), .Y(n791) );
  OAI2B2X1 U2517 ( .A1N(Output2[73]), .A0(n2507), .B0(n2582), .B1(n2508), .Y(
        n792) );
  XOR2X1 U2518 ( .A(n1159), .B(n2583), .Y(Output2[73]) );
  NOR2X1 U2519 ( .A(n246), .B(n2582), .Y(n2583) );
  CLKINVX1 U2520 ( .A(Input2[73]), .Y(n2582) );
  OAI221X1 U2521 ( .A0(n2197), .A1(n2274), .B0(n2203), .B1(n278), .C0(n2584), 
        .Y(n1159) );
  AOI22XL U2522 ( .A0(n262), .A1(n2585), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[75]), .B1(n299), .Y(n2584) );
  MXI2X1 U2523 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[79]), .B(n2586), .S0(
        n307), .Y(n2197) );
  XOR2X1 U2524 ( .A(n2587), .B(n2588), .Y(n2586) );
  XOR2X1 U2525 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[39]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_31_), .Y(n2588) );
  OAI221X1 U2526 ( .A0(n795), .A1(n166), .B0(n1161), .B1(n151), .C0(n2589), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_72_N3) );
  AOI22XL U2527 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_72_), 
        .B0(n234), .B1(Input2[72]), .Y(n2589) );
  CLKINVX1 U2528 ( .A(n796), .Y(n795) );
  OAI2B2X1 U2529 ( .A1N(Input2[72]), .A0(n2508), .B0(n2590), .B1(n2507), .Y(
        n796) );
  CLKINVX1 U2530 ( .A(Output2[72]), .Y(n2590) );
  XOR2X1 U2531 ( .A(n2591), .B(n1161), .Y(Output2[72]) );
  AOI221XL U2532 ( .A0(n2515), .A1(n296), .B0(n2544), .B1(n2293), .C0(n2592), 
        .Y(n1161) );
  AO22X1 U2533 ( .A0(n266), .A1(n2593), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C2[72]), .B1(n292), .Y(n2592) );
  CLKINVX1 U2534 ( .A(n2079), .Y(n2544) );
  MXI2X1 U2535 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[73]), .B(n2594), .S0(
        n307), .Y(n2079) );
  XOR2X1 U2536 ( .A(n2595), .B(n2596), .Y(n2594) );
  XOR2X1 U2537 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[33]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_25_), .Y(n2596) );
  XOR2X1 U2538 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_18_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[72]), .Y(n2515) );
  CLKNAND2X2 U2539 ( .A(Input2[72]), .B(n2288), .Y(n2591) );
  OAI221X1 U2540 ( .A0(n2597), .A1(n2300), .B0(n2598), .B1(n2302), .C0(n2599), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_71_N3) );
  AOI22XL U2541 ( .A0(n186), .A1(n799), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1163), .Y(n2599) );
  OAI2B2X1 U2542 ( .A1N(Output2[71]), .A0(n2600), .B0(n2598), .B1(n2601), .Y(
        n799) );
  XOR2X1 U2543 ( .A(n1163), .B(n2602), .Y(Output2[71]) );
  NOR2X1 U2544 ( .A(n246), .B(n2598), .Y(n2602) );
  OAI221X1 U2545 ( .A0(n2603), .A1(n2273), .B0(n2267), .B1(n2604), .C0(n2605), 
        .Y(n1163) );
  AOI222XL U2546 ( .A0(n290), .A1(n2606), .B0(n2258), .B1(n2607), .C0(n2312), 
        .C1(n2608), .Y(n2605) );
  XOR2X1 U2547 ( .A(n2609), .B(n2610), .Y(n2607) );
  XOR2X1 U2548 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[47]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_37_), .Y(n2610) );
  CLKINVX1 U2549 ( .A(Input2[71]), .Y(n2598) );
  CLKINVX1 U2550 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_71_), .Y(n2597) );
  OAI221X1 U2551 ( .A0(n802), .A1(n165), .B0(n1165), .B1(n151), .C0(n2611), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_70_N3) );
  AOI22XL U2552 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_70_), 
        .B0(n234), .B1(Input2[70]), .Y(n2611) );
  CLKINVX1 U2553 ( .A(n803), .Y(n802) );
  OAI2B2X1 U2554 ( .A1N(Input2[70]), .A0(n2601), .B0(n2612), .B1(n2600), .Y(
        n803) );
  CLKINVX1 U2555 ( .A(Output2[70]), .Y(n2612) );
  XOR2X1 U2556 ( .A(n2613), .B(n1165), .Y(Output2[70]) );
  AOI221XL U2557 ( .A0(n2614), .A1(n2293), .B0(n2615), .B1(n265), .C0(n2616), 
        .Y(n1165) );
  OAI2BB2X1 U2558 ( .B0(n2604), .B1(n284), .A0N(
        Inst_forkAE_CipherInst_RF_S_MID_D2[66]), .A1N(n301), .Y(n2616) );
  CLKINVX1 U2559 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[65]), .Y(n2604) );
  XNOR2X1 U2560 ( .A(n2617), .B(n2618), .Y(n2614) );
  MXI2X1 U2561 ( .A(n2619), .B(n2620), .S0(n307), .Y(n2618) );
  XOR2X1 U2562 ( .A(n2621), .B(n2622), .Y(n2620) );
  XOR2X1 U2563 ( .A(n2623), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[60]), .Y(
        n2621) );
  CLKINVX1 U2564 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[68]), .Y(n2619) );
  OR2X1 U2565 ( .A(n2205), .B(n2083), .Y(n2617) );
  CLKNAND2X2 U2566 ( .A(Input2[70]), .B(n2288), .Y(n2613) );
  OAI221X1 U2567 ( .A0(n2624), .A1(n2300), .B0(n2625), .B1(n2302), .C0(n2626), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_7_N3) );
  AOI22XL U2568 ( .A0(n186), .A1(n1047), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1272), .Y(n2626) );
  AO22X1 U2569 ( .A0(Input2[7]), .A1(n2627), .B0(n1989), .B1(Output2[7]), .Y(
        n1047) );
  XOR2X1 U2570 ( .A(n1272), .B(n2628), .Y(Output2[7]) );
  NOR2X1 U2571 ( .A(n246), .B(n2625), .Y(n2628) );
  OAI221X1 U2572 ( .A0(n2629), .A1(n2273), .B0(n2267), .B1(n2630), .C0(n2631), 
        .Y(n1272) );
  AOI222XL U2573 ( .A0(n291), .A1(n2632), .B0(n2258), .B1(n2633), .C0(n2312), 
        .C1(n2634), .Y(n2631) );
  XOR2X1 U2574 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[104]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[23]), .Y(n2633) );
  CLKINVX1 U2575 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .Y(n2630) );
  CLKINVX1 U2576 ( .A(Input2[7]), .Y(n2625) );
  CLKINVX1 U2577 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_7_), .Y(n2624) );
  OAI221X1 U2578 ( .A0(n806), .A1(n171), .B0(n1166), .B1(n150), .C0(n2635), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_69_N3) );
  AOI22XL U2579 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_69_), 
        .B0(n234), .B1(Input2[69]), .Y(n2635) );
  CLKINVX1 U2580 ( .A(n807), .Y(n806) );
  OAI2B2X1 U2581 ( .A1N(Output2[69]), .A0(n2600), .B0(n2636), .B1(n2601), .Y(
        n807) );
  XNOR2X1 U2582 ( .A(n1166), .B(n2637), .Y(Output2[69]) );
  NOR2X1 U2583 ( .A(n246), .B(n2636), .Y(n2637) );
  CLKINVX1 U2584 ( .A(Input2[69]), .Y(n2636) );
  AOI222XL U2585 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), 
        .B0(n2638), .B1(n2293), .C0(n2639), .C1(n265), .Y(n1166) );
  XNOR2X1 U2586 ( .A(n2640), .B(n2641), .Y(n2638) );
  MXI2X1 U2587 ( .A(n2642), .B(n2643), .S0(n307), .Y(n2641) );
  XOR2X1 U2588 ( .A(n2644), .B(n2645), .Y(n2643) );
  XOR2X1 U2589 ( .A(n2646), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[56]), .Y(
        n2644) );
  CLKNAND2X2 U2590 ( .A(n2647), .B(n2648), .Y(n2640) );
  OAI221X1 U2591 ( .A0(n810), .A1(n177), .B0(n1168), .B1(n150), .C0(n2649), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_68_N3) );
  AOI22XL U2592 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_68_), 
        .B0(n233), .B1(Input2[68]), .Y(n2649) );
  CLKINVX1 U2593 ( .A(n811), .Y(n810) );
  OAI2B2X1 U2594 ( .A1N(Input2[68]), .A0(n2601), .B0(n2650), .B1(n2600), .Y(
        n811) );
  CLKINVX1 U2595 ( .A(Output2[68]), .Y(n2650) );
  XOR2X1 U2596 ( .A(n2651), .B(n1168), .Y(Output2[68]) );
  AOI221XL U2597 ( .A0(n2652), .A1(n296), .B0(n2648), .B1(n2293), .C0(n2653), 
        .Y(n1168) );
  OAI2BB2X1 U2598 ( .B0(n2085), .B1(n284), .A0N(n2654), .A1N(n268), .Y(n2653)
         );
  CLKINVX1 U2599 ( .A(n2209), .Y(n2648) );
  MXI2X1 U2600 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[67]), .B(n2655), .S0(
        n307), .Y(n2209) );
  XOR2X1 U2601 ( .A(n2656), .B(n2657), .Y(n2655) );
  XOR2X1 U2602 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[59]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_35_), .Y(n2657) );
  CLKNAND2X2 U2603 ( .A(Input2[68]), .B(n2288), .Y(n2651) );
  OAI221X1 U2604 ( .A0(n814), .A1(n178), .B0(n2658), .B1(n150), .C0(n2659), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_67_N3) );
  AOI22XL U2605 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_67_), 
        .B0(n233), .B1(Input2[67]), .Y(n2659) );
  CLKINVX1 U2606 ( .A(n1170), .Y(n2658) );
  CLKINVX1 U2607 ( .A(n815), .Y(n814) );
  OAI2B2X1 U2608 ( .A1N(Output2[67]), .A0(n2600), .B0(n2660), .B1(n2601), .Y(
        n815) );
  XOR2X1 U2609 ( .A(n1170), .B(n2661), .Y(Output2[67]) );
  NOR2X1 U2610 ( .A(n246), .B(n2660), .Y(n2661) );
  CLKINVX1 U2611 ( .A(Input2[67]), .Y(n2660) );
  OAI211XL U2612 ( .A0(n2662), .A1(n2273), .B0(n2663), .C0(n2664), .Y(n1170)
         );
  AOI22XL U2613 ( .A0(n2258), .A1(n2665), .B0(n2312), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D2[66]), .Y(n2664) );
  XNOR2X1 U2614 ( .A(n2666), .B(n2667), .Y(n2665) );
  XOR2X1 U2615 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[58]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_34_), .Y(n2667) );
  MXI2X1 U2616 ( .A(n2668), .B(n2669), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[68]), .Y(n2663) );
  OAI21X1 U2617 ( .A0(n2670), .A1(n279), .B0(n2267), .Y(n2669) );
  NOR2X1 U2618 ( .A(n2085), .B(n2207), .Y(n2670) );
  NOR3X1 U2619 ( .A(n2207), .B(n276), .C(n2085), .Y(n2668) );
  CLKINVX1 U2620 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[68]), .Y(n2085) );
  CLKINVX1 U2621 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), .Y(n2207) );
  OAI221X1 U2622 ( .A0(n818), .A1(n179), .B0(n1171), .B1(n150), .C0(n2671), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_66_N3) );
  AOI22XL U2623 ( .A0(n206), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_66_), 
        .B0(n233), .B1(Input2[66]), .Y(n2671) );
  CLKINVX1 U2624 ( .A(n819), .Y(n818) );
  OAI2B2X1 U2625 ( .A1N(Output2[66]), .A0(n2600), .B0(n2672), .B1(n2601), .Y(
        n819) );
  XNOR2X1 U2626 ( .A(n1171), .B(n2673), .Y(Output2[66]) );
  NOR2X1 U2627 ( .A(n246), .B(n2672), .Y(n2673) );
  CLKINVX1 U2628 ( .A(Input2[66]), .Y(n2672) );
  AOI221XL U2629 ( .A0(n2674), .A1(n2293), .B0(n2675), .B1(n265), .C0(n2676), 
        .Y(n1171) );
  MX2X1 U2630 ( .A(n2677), .B(n2678), .S0(n2642), .Y(n2676) );
  CLKINVX1 U2631 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[64]), .Y(n2642) );
  NOR3X1 U2632 ( .A(n277), .B(n2088), .C(n2211), .Y(n2678) );
  OAI21X1 U2633 ( .A0(n2679), .A1(n279), .B0(n2267), .Y(n2677) );
  NOR2X1 U2634 ( .A(n2088), .B(n2211), .Y(n2679) );
  CLKINVX1 U2635 ( .A(n2083), .Y(n2674) );
  MXI2X1 U2636 ( .A(n2652), .B(n2680), .S0(n307), .Y(n2083) );
  XOR2X1 U2637 ( .A(n2681), .B(n2682), .Y(n2680) );
  XOR2X1 U2638 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[42]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_), .Y(n2682) );
  XOR2X1 U2639 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_17_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[68]), .Y(n2652) );
  OAI221X1 U2640 ( .A0(n822), .A1(n179), .B0(n2683), .B1(n150), .C0(n2684), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_65_N3) );
  AOI22XL U2641 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_65_), 
        .B0(n233), .B1(Input2[65]), .Y(n2684) );
  CLKINVX1 U2642 ( .A(n1173), .Y(n2683) );
  CLKINVX1 U2643 ( .A(n823), .Y(n822) );
  OAI2B2X1 U2644 ( .A1N(Output2[65]), .A0(n2600), .B0(n2685), .B1(n2601), .Y(
        n823) );
  XOR2X1 U2645 ( .A(n1173), .B(n2686), .Y(Output2[65]) );
  NOR2X1 U2646 ( .A(n246), .B(n2685), .Y(n2686) );
  CLKINVX1 U2647 ( .A(Input2[65]), .Y(n2685) );
  OAI221X1 U2648 ( .A0(n2205), .A1(n2274), .B0(n2211), .B1(n278), .C0(n2687), 
        .Y(n1173) );
  AOI22XL U2649 ( .A0(n261), .A1(n2688), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[67]), .B1(n300), .Y(n2687) );
  MXI2X1 U2650 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), .B(n2689), .S0(
        n307), .Y(n2205) );
  XOR2X1 U2651 ( .A(n2690), .B(n2691), .Y(n2689) );
  XOR2X1 U2652 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[63]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_39_), .Y(n2691) );
  OAI221X1 U2653 ( .A0(n826), .A1(n179), .B0(n1175), .B1(n150), .C0(n2692), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_64_N3) );
  AOI22XL U2654 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_64_), 
        .B0(n233), .B1(Input2[64]), .Y(n2692) );
  CLKINVX1 U2655 ( .A(n827), .Y(n826) );
  OAI2B2X1 U2656 ( .A1N(Input2[64]), .A0(n2601), .B0(n2693), .B1(n2600), .Y(
        n827) );
  CLKINVX1 U2657 ( .A(Output2[64]), .Y(n2693) );
  XOR2X1 U2658 ( .A(n2694), .B(n1175), .Y(Output2[64]) );
  AOI221XL U2659 ( .A0(n2608), .A1(n296), .B0(n2647), .B1(n2293), .C0(n2695), 
        .Y(n1175) );
  AO22X1 U2660 ( .A0(n266), .A1(n2696), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C2[64]), .B1(n292), .Y(n2695) );
  CLKINVX1 U2661 ( .A(n2086), .Y(n2647) );
  MXI2X1 U2662 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[65]), .B(n2697), .S0(
        n307), .Y(n2086) );
  XOR2X1 U2663 ( .A(n2698), .B(n2699), .Y(n2697) );
  XOR2X1 U2664 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[57]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_33_), .Y(n2699) );
  XOR2X1 U2665 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_16_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[64]), .Y(n2608) );
  CLKNAND2X2 U2666 ( .A(Input2[64]), .B(n2288), .Y(n2694) );
  OAI221X1 U2667 ( .A0(n2700), .A1(n2300), .B0(n2701), .B1(n2302), .C0(n2702), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_63_N3) );
  AOI22XL U2668 ( .A0(n186), .A1(n830), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1177), .Y(n2702) );
  OAI2B2X1 U2669 ( .A1N(Output2[63]), .A0(n2703), .B0(n2701), .B1(n2704), .Y(
        n830) );
  XOR2X1 U2670 ( .A(n1177), .B(n2705), .Y(Output2[63]) );
  NOR2X1 U2671 ( .A(n246), .B(n2701), .Y(n2705) );
  OAI221X1 U2672 ( .A0(n2095), .A1(n277), .B0(n2267), .B1(n2706), .C0(n2707), 
        .Y(n1177) );
  AOI222XL U2673 ( .A0(n2258), .A1(n2416), .B0(n260), .B1(n2708), .C0(n2312), 
        .C1(n2709), .Y(n2707) );
  XOR2X1 U2674 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_39_), .B(n2710), 
        .Y(n2708) );
  XOR2X1 U2675 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[64]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[63]), .Y(n2710) );
  XOR2X1 U2676 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[23]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[72]), .Y(n2416) );
  CLKINVX1 U2677 ( .A(Input2[63]), .Y(n2701) );
  CLKINVX1 U2678 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_63_), .Y(n2700) );
  OAI221X1 U2679 ( .A0(n833), .A1(n179), .B0(n1178), .B1(n150), .C0(n2711), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_62_N3) );
  AOI22XL U2680 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_62_), 
        .B0(n233), .B1(Input2[62]), .Y(n2711) );
  CLKINVX1 U2681 ( .A(n834), .Y(n833) );
  OAI2B2X1 U2682 ( .A1N(Output2[62]), .A0(n2703), .B0(n2712), .B1(n2704), .Y(
        n834) );
  CLKINVX1 U2683 ( .A(Input2[62]), .Y(n2712) );
  XOR2X1 U2684 ( .A(n2713), .B(n1178), .Y(Output2[62]) );
  CLKINVX1 U2685 ( .A(n2714), .Y(n1178) );
  OAI211XL U2686 ( .A0(n285), .A1(n2706), .B0(n2715), .C0(n2716), .Y(n2714) );
  AOI22XL U2687 ( .A0(n262), .A1(n2717), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[58]), .B1(n300), .Y(n2716) );
  XOR2X1 U2688 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_), .B(n2718), 
        .Y(n2717) );
  XOR2X1 U2689 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[68]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[44]), .Y(n2718) );
  MXI2X1 U2690 ( .A(n2719), .B(n2720), .S0(n2721), .Y(n2715) );
  NOR2X1 U2691 ( .A(n2090), .B(n2213), .Y(n2721) );
  OAI22X1 U2692 ( .A0(n2722), .A1(n2429), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[60]), .B1(n2255), .Y(n2720) );
  OAI2BB2X1 U2693 ( .B0(n2255), .B1(n2723), .A0N(n2429), .A1N(n2258), .Y(n2719) );
  XNOR2X1 U2694 ( .A(n2724), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[76]), .Y(
        n2429) );
  CLKNAND2X2 U2695 ( .A(Input2[62]), .B(n2288), .Y(n2713) );
  OAI221X1 U2696 ( .A0(n837), .A1(n179), .B0(n1179), .B1(n150), .C0(n2725), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_61_N3) );
  AOI22XL U2697 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_61_), 
        .B0(n233), .B1(Input2[61]), .Y(n2725) );
  CLKINVX1 U2698 ( .A(n838), .Y(n837) );
  OAI2B2X1 U2699 ( .A1N(Output2[61]), .A0(n2703), .B0(n2726), .B1(n2704), .Y(
        n838) );
  CLKINVX1 U2700 ( .A(Input2[61]), .Y(n2726) );
  XOR2X1 U2701 ( .A(n2727), .B(n1179), .Y(Output2[61]) );
  CLKINVX1 U2702 ( .A(n2728), .Y(n1179) );
  OAI221X1 U2703 ( .A0(n2729), .A1(n2273), .B0(n2730), .B1(n2215), .C0(n2731), 
        .Y(n2728) );
  MXI2X1 U2704 ( .A(n2732), .B(n2733), .S0(n2734), .Y(n2731) );
  NOR2X1 U2705 ( .A(n2216), .B(n2093), .Y(n2734) );
  OAI22X1 U2706 ( .A0(n2722), .A1(n2441), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[56]), .B1(n2255), .Y(n2733) );
  OAI2BB2X1 U2707 ( .B0(n2255), .B1(n2735), .A0N(n2441), .A1N(n2258), .Y(n2732) );
  XNOR2X1 U2708 ( .A(n2539), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[8]), .Y(
        n2441) );
  CLKINVX1 U2709 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[72]), .Y(n2539) );
  XOR2X1 U2710 ( .A(n2736), .B(n2737), .Y(n2729) );
  XOR2X1 U2711 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[64]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[40]), .Y(n2737) );
  CLKNAND2X2 U2712 ( .A(Input2[61]), .B(n2288), .Y(n2727) );
  OAI221X1 U2713 ( .A0(n841), .A1(n179), .B0(n2738), .B1(n150), .C0(n2739), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_60_N3) );
  AOI22XL U2714 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_60_), 
        .B0(n233), .B1(Input2[60]), .Y(n2739) );
  CLKINVX1 U2715 ( .A(n1181), .Y(n2738) );
  CLKINVX1 U2716 ( .A(n842), .Y(n841) );
  OAI2B2X1 U2717 ( .A1N(Output2[60]), .A0(n2703), .B0(n2740), .B1(n2704), .Y(
        n842) );
  XOR2X1 U2718 ( .A(n1181), .B(n2741), .Y(Output2[60]) );
  NOR2X1 U2719 ( .A(n246), .B(n2740), .Y(n2741) );
  CLKINVX1 U2720 ( .A(Input2[60]), .Y(n2740) );
  OAI221X1 U2721 ( .A0(n2216), .A1(n2274), .B0(n285), .B1(n2092), .C0(n2742), 
        .Y(n1181) );
  AOI22XL U2722 ( .A0(n261), .A1(n2743), .B0(n294), .B1(n2744), .Y(n2742) );
  XOR2X1 U2723 ( .A(n2745), .B(n2746), .Y(n2743) );
  XOR2X1 U2724 ( .A(n2623), .B(n2211), .Y(n2746) );
  XNOR2X1 U2725 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_17_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[67]), .Y(n2211) );
  MXI2X1 U2726 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[59]), .B(n2452), .S0(
        n308), .Y(n2216) );
  XOR2X1 U2727 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[11]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[75]), .Y(n2452) );
  OAI221X1 U2728 ( .A0(n1050), .A1(n179), .B0(n1273), .B1(n150), .C0(n2747), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_6_N3) );
  AOI22XL U2729 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_6_), 
        .B0(n233), .B1(Input2[6]), .Y(n2747) );
  AOI22XL U2730 ( .A0(Input2[6]), .A1(n2627), .B0(n1989), .B1(Output2[6]), .Y(
        n1050) );
  XOR2X1 U2731 ( .A(n2748), .B(n1273), .Y(Output2[6]) );
  CLKINVX1 U2732 ( .A(n2749), .Y(n1273) );
  OAI221X1 U2733 ( .A0(n2750), .A1(n2274), .B0(n2751), .B1(n2273), .C0(n2752), 
        .Y(n2749) );
  AOI22XL U2734 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[2]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .B1(n292), .Y(n2752) );
  XOR2X1 U2735 ( .A(n2753), .B(n2754), .Y(n2750) );
  MXI2X1 U2736 ( .A(n2755), .B(n2756), .S0(n308), .Y(n2754) );
  XOR2X1 U2737 ( .A(n2757), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[12]), .Y(
        n2756) );
  OR2X1 U2738 ( .A(n2141), .B(n2022), .Y(n2753) );
  CLKNAND2X2 U2739 ( .A(Input2[6]), .B(n2288), .Y(n2748) );
  OAI221X1 U2740 ( .A0(n845), .A1(n179), .B0(n2758), .B1(n150), .C0(n2759), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_59_N3) );
  AOI22XL U2741 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_59_), 
        .B0(n233), .B1(Input2[59]), .Y(n2759) );
  CLKINVX1 U2742 ( .A(n1183), .Y(n2758) );
  CLKINVX1 U2743 ( .A(n846), .Y(n845) );
  OAI2B2X1 U2744 ( .A1N(Output2[59]), .A0(n2703), .B0(n2760), .B1(n2704), .Y(
        n846) );
  XOR2X1 U2745 ( .A(n1183), .B(n2761), .Y(Output2[59]) );
  NOR2X1 U2746 ( .A(n246), .B(n2760), .Y(n2761) );
  CLKINVX1 U2747 ( .A(Input2[59]), .Y(n2760) );
  OAI211XL U2748 ( .A0(n2462), .A1(n2722), .B0(n2762), .C0(n2763), .Y(n1183)
         );
  AOI22XL U2749 ( .A0(n262), .A1(n2764), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[58]), .B1(n2312), .Y(n2763) );
  XOR2X1 U2750 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_35_), .B(n2765), 
        .Y(n2764) );
  XOR2X1 U2751 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[65]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[41]), .Y(n2765) );
  MXI2X1 U2752 ( .A(n2766), .B(n2767), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[60]), .Y(n2762) );
  OAI21X1 U2753 ( .A0(n2768), .A1(n279), .B0(n2267), .Y(n2767) );
  NOR2X1 U2754 ( .A(n2215), .B(n2092), .Y(n2768) );
  NOR3X1 U2755 ( .A(n2092), .B(n2215), .C(n278), .Y(n2766) );
  XNOR2X1 U2756 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[74]), .Y(n2462) );
  OAI221X1 U2757 ( .A0(n849), .A1(n179), .B0(n2769), .B1(n150), .C0(n2770), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_58_N3) );
  AOI22XL U2758 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_58_), 
        .B0(n233), .B1(Input2[58]), .Y(n2770) );
  CLKINVX1 U2759 ( .A(n1185), .Y(n2769) );
  CLKINVX1 U2760 ( .A(n850), .Y(n849) );
  OAI2B2X1 U2761 ( .A1N(Output2[58]), .A0(n2703), .B0(n2771), .B1(n2704), .Y(
        n850) );
  XOR2X1 U2762 ( .A(n1185), .B(n2772), .Y(Output2[58]) );
  NOR2X1 U2763 ( .A(n246), .B(n2771), .Y(n2772) );
  CLKINVX1 U2764 ( .A(Input2[58]), .Y(n2771) );
  OAI221X1 U2765 ( .A0(n2773), .A1(n2273), .B0(n2090), .B1(n2274), .C0(n2774), 
        .Y(n1185) );
  MXI2X1 U2766 ( .A(n2775), .B(n2776), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[56]), .Y(n2774) );
  OAI21X1 U2767 ( .A0(n2777), .A1(n279), .B0(n2267), .Y(n2776) );
  NOR2X1 U2768 ( .A(n2095), .B(n2218), .Y(n2777) );
  NOR3X1 U2769 ( .A(n275), .B(n2095), .C(n2218), .Y(n2775) );
  MXI2X1 U2770 ( .A(n2744), .B(n2477), .S0(n308), .Y(n2090) );
  XOR2X1 U2771 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[76]), .Y(n2477) );
  XOR2X1 U2772 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_15_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[42]), .Y(n2744) );
  XOR2X1 U2773 ( .A(n2778), .B(n2779), .Y(n2773) );
  XOR2X1 U2774 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[68]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[58]), .Y(n2779) );
  OAI221X1 U2775 ( .A0(n853), .A1(n179), .B0(n1186), .B1(n150), .C0(n2780), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_57_N3) );
  AOI22XL U2776 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_57_), 
        .B0(n233), .B1(Input2[57]), .Y(n2780) );
  CLKINVX1 U2777 ( .A(n854), .Y(n853) );
  OAI2B2X1 U2778 ( .A1N(Output2[57]), .A0(n2703), .B0(n2781), .B1(n2704), .Y(
        n854) );
  CLKINVX1 U2779 ( .A(Input2[57]), .Y(n2781) );
  XOR2X1 U2780 ( .A(n2782), .B(n1186), .Y(Output2[57]) );
  CLKINVX1 U2781 ( .A(n2783), .Y(n1186) );
  OAI221X1 U2782 ( .A0(n2784), .A1(n2273), .B0(n2213), .B1(n2274), .C0(n2785), 
        .Y(n2783) );
  AOI22XL U2783 ( .A0(n291), .A1(n2786), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[59]), .B1(n300), .Y(n2785) );
  MXI2X1 U2784 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[63]), .B(n2486), .S0(
        n308), .Y(n2213) );
  XOR2X1 U2785 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[79]), .Y(n2486) );
  XOR2X1 U2786 ( .A(n2787), .B(n2788), .Y(n2784) );
  XOR2X1 U2787 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[47]), .Y(n2788) );
  CLKNAND2X2 U2788 ( .A(Input2[57]), .B(n2288), .Y(n2782) );
  OAI221X1 U2789 ( .A0(n857), .A1(n179), .B0(n2789), .B1(n150), .C0(n2790), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_56_N3) );
  AOI22XL U2790 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_56_), 
        .B0(n233), .B1(Input2[56]), .Y(n2790) );
  CLKINVX1 U2791 ( .A(n1188), .Y(n2789) );
  CLKINVX1 U2792 ( .A(n858), .Y(n857) );
  OAI2B2X1 U2793 ( .A1N(Output2[56]), .A0(n2703), .B0(n2791), .B1(n2704), .Y(
        n858) );
  XOR2X1 U2794 ( .A(n1188), .B(n2792), .Y(Output2[56]) );
  NOR2X1 U2795 ( .A(n246), .B(n2791), .Y(n2792) );
  CLKINVX1 U2796 ( .A(Input2[56]), .Y(n2791) );
  OAI221X1 U2797 ( .A0(n2093), .A1(n2274), .B0(n2266), .B1(n2793), .C0(n2794), 
        .Y(n1188) );
  AOI22XL U2798 ( .A0(n262), .A1(n2795), .B0(n294), .B1(n2709), .Y(n2794) );
  XNOR2X1 U2799 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_14_), .B(n2793), .Y(
        n2709) );
  XOR2X1 U2800 ( .A(n2796), .B(n2797), .Y(n2795) );
  XOR2X1 U2801 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_32_), .B(n2606), 
        .Y(n2797) );
  CLKINVX1 U2802 ( .A(n2088), .Y(n2606) );
  XNOR2X1 U2803 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_16_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[66]), .Y(n2088) );
  CLKINVX1 U2804 ( .A(n2109), .Y(n2796) );
  CLKINVX1 U2805 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[47]), .Y(n2793) );
  MXI2X1 U2806 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[57]), .B(n2494), .S0(
        n308), .Y(n2093) );
  XOR2X1 U2807 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[73]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .Y(n2494) );
  OAI221X1 U2808 ( .A0(n2798), .A1(n2300), .B0(n2799), .B1(n2302), .C0(n2800), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_55_N3) );
  AOI22XL U2809 ( .A0(n186), .A1(n861), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1190), .Y(n2800) );
  OAI2B2X1 U2810 ( .A1N(Output2[55]), .A0(n2801), .B0(n2799), .B1(n2802), .Y(
        n861) );
  XOR2X1 U2811 ( .A(n1190), .B(n2803), .Y(Output2[55]) );
  NOR2X1 U2812 ( .A(n246), .B(n2799), .Y(n2803) );
  OAI221X1 U2813 ( .A0(n2102), .A1(n277), .B0(n2267), .B1(n2804), .C0(n2805), 
        .Y(n1190) );
  AOI222XL U2814 ( .A0(n2258), .A1(n2516), .B0(n260), .B1(n2806), .C0(n2312), 
        .C1(n2807), .Y(n2805) );
  XOR2X1 U2815 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_47_), .B(n2808), 
        .Y(n2806) );
  XOR2X1 U2816 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[88]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[55]), .Y(n2808) );
  XOR2X1 U2817 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[64]), .Y(n2516) );
  CLKINVX1 U2818 ( .A(Input2[55]), .Y(n2799) );
  CLKINVX1 U2819 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_55_), .Y(n2798) );
  OAI221X1 U2820 ( .A0(n864), .A1(n179), .B0(n1191), .B1(n150), .C0(n2809), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_54_N3) );
  AOI22XL U2821 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_54_), 
        .B0(n232), .B1(Input2[54]), .Y(n2809) );
  CLKINVX1 U2822 ( .A(n865), .Y(n864) );
  OAI2B2X1 U2823 ( .A1N(Output2[54]), .A0(n2801), .B0(n2810), .B1(n2802), .Y(
        n865) );
  CLKINVX1 U2824 ( .A(Input2[54]), .Y(n2810) );
  XOR2X1 U2825 ( .A(n2811), .B(n1191), .Y(Output2[54]) );
  CLKINVX1 U2826 ( .A(n2812), .Y(n1191) );
  OAI211XL U2827 ( .A0(n285), .A1(n2804), .B0(n2813), .C0(n2814), .Y(n2812) );
  AOI22XL U2828 ( .A0(n263), .A1(n2815), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[50]), .B1(n299), .Y(n2814) );
  XOR2X1 U2829 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_), .B(n2816), 
        .Y(n2815) );
  XOR2X1 U2830 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[92]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[36]), .Y(n2816) );
  MXI2X1 U2831 ( .A(n2817), .B(n2818), .S0(n2819), .Y(n2813) );
  NOR2X1 U2832 ( .A(n2097), .B(n2220), .Y(n2819) );
  OAI22X1 U2833 ( .A0(n2722), .A1(n2530), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .B1(n2255), .Y(n2818) );
  AO22X1 U2834 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .A1(n2312), .B0(
        n2530), .B1(n2258), .Y(n2817) );
  XNOR2X1 U2835 ( .A(n2755), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[68]), .Y(
        n2530) );
  CLKINVX1 U2836 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[4]), .Y(n2755) );
  CLKNAND2X2 U2837 ( .A(Input2[54]), .B(n2288), .Y(n2811) );
  OAI221X1 U2838 ( .A0(n868), .A1(n179), .B0(n1192), .B1(n150), .C0(n2820), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_53_N3) );
  AOI22XL U2839 ( .A0(n205), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_53_), 
        .B0(n232), .B1(Input2[53]), .Y(n2820) );
  CLKINVX1 U2840 ( .A(n869), .Y(n868) );
  OAI2B2X1 U2841 ( .A1N(Output2[53]), .A0(n2801), .B0(n2821), .B1(n2802), .Y(
        n869) );
  CLKINVX1 U2842 ( .A(Input2[53]), .Y(n2821) );
  XOR2X1 U2843 ( .A(n2822), .B(n1192), .Y(Output2[53]) );
  CLKINVX1 U2844 ( .A(n2823), .Y(n1192) );
  OAI221X1 U2845 ( .A0(n2824), .A1(n2273), .B0(n2730), .B1(n2222), .C0(n2825), 
        .Y(n2823) );
  MXI2X1 U2846 ( .A(n2826), .B(n2827), .S0(n2828), .Y(n2825) );
  NOR2X1 U2847 ( .A(n2223), .B(n2100), .Y(n2828) );
  OAI22X1 U2848 ( .A0(n2722), .A1(n2542), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .B1(n2255), .Y(n2827) );
  AO22X1 U2849 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .A1(n2312), .B0(
        n2542), .B1(n2258), .Y(n2826) );
  XNOR2X1 U2850 ( .A(n2829), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[64]), .Y(
        n2542) );
  XOR2X1 U2851 ( .A(n2830), .B(n2831), .Y(n2824) );
  XOR2X1 U2852 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[88]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[32]), .Y(n2831) );
  CLKNAND2X2 U2853 ( .A(Input2[53]), .B(n2288), .Y(n2822) );
  OAI221X1 U2854 ( .A0(n872), .A1(n178), .B0(n2832), .B1(n149), .C0(n2833), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_52_N3) );
  AOI22XL U2855 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_52_), 
        .B0(n232), .B1(Input2[52]), .Y(n2833) );
  CLKINVX1 U2856 ( .A(n1194), .Y(n2832) );
  CLKINVX1 U2857 ( .A(n873), .Y(n872) );
  OAI2B2X1 U2858 ( .A1N(Output2[52]), .A0(n2801), .B0(n2834), .B1(n2802), .Y(
        n873) );
  XOR2X1 U2859 ( .A(n1194), .B(n2835), .Y(Output2[52]) );
  NOR2X1 U2860 ( .A(n247), .B(n2834), .Y(n2835) );
  CLKINVX1 U2861 ( .A(Input2[52]), .Y(n2834) );
  OAI221X1 U2862 ( .A0(n2223), .A1(n2274), .B0(n279), .B1(n2099), .C0(n2836), 
        .Y(n1194) );
  AOI22XL U2863 ( .A0(n263), .A1(n2837), .B0(n295), .B1(n2838), .Y(n2836) );
  XOR2X1 U2864 ( .A(n2839), .B(n2840), .Y(n2837) );
  XOR2X1 U2865 ( .A(n2328), .B(n2187), .Y(n2840) );
  XNOR2X1 U2866 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_23_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[91]), .Y(n2187) );
  MXI2X1 U2867 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[51]), .B(n2553), .S0(
        n308), .Y(n2223) );
  XOR2X1 U2868 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[3]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[67]), .Y(n2553) );
  OAI221X1 U2869 ( .A0(n876), .A1(n178), .B0(n2841), .B1(n149), .C0(n2842), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_51_N3) );
  AOI22XL U2870 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_51_), 
        .B0(n232), .B1(Input2[51]), .Y(n2842) );
  CLKINVX1 U2871 ( .A(n1196), .Y(n2841) );
  CLKINVX1 U2872 ( .A(n877), .Y(n876) );
  OAI2B2X1 U2873 ( .A1N(Output2[51]), .A0(n2801), .B0(n2843), .B1(n2802), .Y(
        n877) );
  XOR2X1 U2874 ( .A(n1196), .B(n2844), .Y(Output2[51]) );
  NOR2X1 U2875 ( .A(n247), .B(n2843), .Y(n2844) );
  CLKINVX1 U2876 ( .A(Input2[51]), .Y(n2843) );
  OAI211XL U2877 ( .A0(n2563), .A1(n2722), .B0(n2845), .C0(n2846), .Y(n1196)
         );
  AOI22XL U2878 ( .A0(n263), .A1(n2847), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[50]), .B1(n2312), .Y(n2846) );
  XOR2X1 U2879 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_43_), .B(n2848), 
        .Y(n2847) );
  XOR2X1 U2880 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[33]), .Y(n2848) );
  MXI2X1 U2881 ( .A(n2849), .B(n2850), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .Y(n2845) );
  OAI21X1 U2882 ( .A0(n2851), .A1(n280), .B0(n2267), .Y(n2850) );
  NOR2X1 U2883 ( .A(n2099), .B(n2222), .Y(n2851) );
  NOR3X1 U2884 ( .A(n2222), .B(n276), .C(n2099), .Y(n2849) );
  XNOR2X1 U2885 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[2]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[66]), .Y(n2563) );
  OAI221X1 U2886 ( .A0(n880), .A1(n178), .B0(n2852), .B1(n149), .C0(n2853), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_50_N3) );
  AOI22XL U2887 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_50_), 
        .B0(n232), .B1(Input2[50]), .Y(n2853) );
  CLKINVX1 U2888 ( .A(n1198), .Y(n2852) );
  CLKINVX1 U2889 ( .A(n881), .Y(n880) );
  OAI2B2X1 U2890 ( .A1N(Output2[50]), .A0(n2801), .B0(n2854), .B1(n2802), .Y(
        n881) );
  XOR2X1 U2891 ( .A(n1198), .B(n2855), .Y(Output2[50]) );
  NOR2X1 U2892 ( .A(n247), .B(n2854), .Y(n2855) );
  CLKINVX1 U2893 ( .A(Input2[50]), .Y(n2854) );
  OAI221X1 U2894 ( .A0(n2856), .A1(n2273), .B0(n2097), .B1(n2274), .C0(n2857), 
        .Y(n1198) );
  MXI2X1 U2895 ( .A(n2858), .B(n2859), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .Y(n2857) );
  OAI21X1 U2896 ( .A0(n2860), .A1(n279), .B0(n2267), .Y(n2859) );
  NOR2X1 U2897 ( .A(n2102), .B(n2225), .Y(n2860) );
  NOR3X1 U2898 ( .A(n275), .B(n2102), .C(n2225), .Y(n2858) );
  MXI2X1 U2899 ( .A(n2838), .B(n2578), .S0(n308), .Y(n2097) );
  XOR2X1 U2900 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[68]), .Y(n2578) );
  XOR2X1 U2901 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_13_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[34]), .Y(n2838) );
  XOR2X1 U2902 ( .A(n2861), .B(n2862), .Y(n2856) );
  XOR2X1 U2903 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[92]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[50]), .Y(n2862) );
  OAI221X1 U2904 ( .A0(n1053), .A1(n178), .B0(n2863), .B1(n149), .C0(n2864), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_5_N3) );
  AOI22XL U2905 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_5_), 
        .B0(n232), .B1(Input2[5]), .Y(n2864) );
  CLKINVX1 U2906 ( .A(n1275), .Y(n2863) );
  AOI22XL U2907 ( .A0(n1989), .A1(Output2[5]), .B0(Input2[5]), .B1(n2627), .Y(
        n1053) );
  XOR2X1 U2908 ( .A(n1275), .B(n2865), .Y(Output2[5]) );
  NOR2BX1 U2909 ( .AN(Input2[5]), .B(n255), .Y(n2865) );
  OAI222X1 U2910 ( .A0(n2730), .A1(n2143), .B0(n2866), .B1(n2274), .C0(n2867), 
        .C1(n2273), .Y(n1275) );
  XOR2X1 U2911 ( .A(n2868), .B(n2869), .Y(n2866) );
  MXI2X1 U2912 ( .A(n2829), .B(n2870), .S0(n308), .Y(n2869) );
  XOR2X1 U2913 ( .A(n2871), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[8]), .Y(
        n2870) );
  CLKNAND2X2 U2914 ( .A(n2872), .B(n2873), .Y(n2868) );
  OAI221X1 U2915 ( .A0(n884), .A1(n178), .B0(n1199), .B1(n149), .C0(n2874), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_49_N3) );
  AOI22XL U2916 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_49_), 
        .B0(n232), .B1(Input2[49]), .Y(n2874) );
  CLKINVX1 U2917 ( .A(n885), .Y(n884) );
  OAI2B2X1 U2918 ( .A1N(Output2[49]), .A0(n2801), .B0(n2875), .B1(n2802), .Y(
        n885) );
  CLKINVX1 U2919 ( .A(Input2[49]), .Y(n2875) );
  XOR2X1 U2920 ( .A(n2876), .B(n1199), .Y(Output2[49]) );
  CLKINVX1 U2921 ( .A(n2877), .Y(n1199) );
  OAI221X1 U2922 ( .A0(n2878), .A1(n2273), .B0(n2220), .B1(n2274), .C0(n2879), 
        .Y(n2877) );
  AOI2BB2X1 U2923 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[51]), .B1(n294), 
        .A0N(n285), .A1N(n2225), .Y(n2879) );
  MXI2X1 U2924 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[55]), .B(n2587), .S0(
        n308), .Y(n2220) );
  XOR2X1 U2925 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[7]), .Y(n2587) );
  XOR2X1 U2926 ( .A(n2880), .B(n2881), .Y(n2878) );
  XOR2X1 U2927 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[95]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[39]), .Y(n2881) );
  CLKNAND2X2 U2928 ( .A(Input2[49]), .B(n2288), .Y(n2876) );
  OAI221X1 U2929 ( .A0(n888), .A1(n178), .B0(n2882), .B1(n149), .C0(n2883), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_48_N3) );
  AOI22XL U2930 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_48_), 
        .B0(n232), .B1(Input2[48]), .Y(n2883) );
  CLKINVX1 U2931 ( .A(n1201), .Y(n2882) );
  CLKINVX1 U2932 ( .A(n889), .Y(n888) );
  OAI2B2X1 U2933 ( .A1N(Output2[48]), .A0(n2801), .B0(n2884), .B1(n2802), .Y(
        n889) );
  XOR2X1 U2934 ( .A(n1201), .B(n2885), .Y(Output2[48]) );
  NOR2X1 U2935 ( .A(n247), .B(n2884), .Y(n2885) );
  CLKINVX1 U2936 ( .A(Input2[48]), .Y(n2884) );
  OAI221X1 U2937 ( .A0(n2100), .A1(n2274), .B0(n280), .B1(n2886), .C0(n2887), 
        .Y(n1201) );
  AOI22XL U2938 ( .A0(n262), .A1(n2888), .B0(n294), .B1(n2807), .Y(n2887) );
  XNOR2X1 U2939 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_12_), .B(n2886), .Y(
        n2807) );
  XOR2X1 U2940 ( .A(n2889), .B(n2890), .Y(n2888) );
  XOR2X1 U2941 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_40_), .B(n2310), 
        .Y(n2890) );
  CLKINVX1 U2942 ( .A(n2067), .Y(n2310) );
  XNOR2X1 U2943 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_22_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[90]), .Y(n2067) );
  CLKINVX1 U2944 ( .A(n2116), .Y(n2889) );
  CLKINVX1 U2945 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[39]), .Y(n2886) );
  MXI2X1 U2946 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[49]), .B(n2595), .S0(
        n308), .Y(n2100) );
  XOR2X1 U2947 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[65]), .Y(n2595) );
  OAI221X1 U2948 ( .A0(n2891), .A1(n2300), .B0(n2892), .B1(n2302), .C0(n2893), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_47_N3) );
  AOI22XL U2949 ( .A0(n186), .A1(n892), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1203), .Y(n2893) );
  OAI2B2X1 U2950 ( .A1N(Output2[47]), .A0(n2894), .B0(n2892), .B1(n2895), .Y(
        n892) );
  XOR2X1 U2951 ( .A(n1203), .B(n2896), .Y(Output2[47]) );
  NOR2X1 U2952 ( .A(n247), .B(n2892), .Y(n2896) );
  OAI221X1 U2953 ( .A0(n2109), .A1(n277), .B0(n2267), .B1(n2897), .C0(n2898), 
        .Y(n1203) );
  AOI222XL U2954 ( .A0(n2258), .A1(n2609), .B0(n260), .B1(n2899), .C0(n2312), 
        .C1(n2900), .Y(n2898) );
  XOR2X1 U2955 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_15_), .B(n2901), 
        .Y(n2899) );
  XOR2X1 U2956 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[80]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[47]), .Y(n2901) );
  XOR2X1 U2957 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[88]), .Y(n2609) );
  CLKINVX1 U2958 ( .A(Input2[47]), .Y(n2892) );
  CLKINVX1 U2959 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_47_), .Y(n2891) );
  OAI221X1 U2960 ( .A0(n895), .A1(n178), .B0(n1204), .B1(n149), .C0(n2902), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_46_N3) );
  AOI22XL U2961 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_46_), 
        .B0(n232), .B1(Input2[46]), .Y(n2902) );
  CLKINVX1 U2962 ( .A(n896), .Y(n895) );
  OAI2B2X1 U2963 ( .A1N(Output2[46]), .A0(n2894), .B0(n2903), .B1(n2895), .Y(
        n896) );
  CLKINVX1 U2964 ( .A(Input2[46]), .Y(n2903) );
  XOR2X1 U2965 ( .A(n2904), .B(n1204), .Y(Output2[46]) );
  CLKINVX1 U2966 ( .A(n2905), .Y(n1204) );
  OAI211XL U2967 ( .A0(n285), .A1(n2897), .B0(n2906), .C0(n2907), .Y(n2905) );
  AOI22XL U2968 ( .A0(n263), .A1(n2908), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[42]), .B1(n300), .Y(n2907) );
  XOR2X1 U2969 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_14_), .B(n2909), 
        .Y(n2908) );
  XOR2X1 U2970 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[84]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[60]), .Y(n2909) );
  MXI2X1 U2971 ( .A(n2910), .B(n2911), .S0(n2912), .Y(n2906) );
  NOR2X1 U2972 ( .A(n2104), .B(n2227), .Y(n2912) );
  OAI22X1 U2973 ( .A0(n2722), .A1(n2622), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[44]), .B1(n2255), .Y(n2911) );
  OAI2BB2X1 U2974 ( .B0(n2255), .B1(n2913), .A0N(n2622), .A1N(n2258), .Y(n2910) );
  XNOR2X1 U2975 ( .A(n2914), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[92]), .Y(
        n2622) );
  CLKNAND2X2 U2976 ( .A(Input2[46]), .B(n2288), .Y(n2904) );
  OAI221X1 U2977 ( .A0(n899), .A1(n178), .B0(n1205), .B1(n149), .C0(n2915), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_45_N3) );
  AOI22XL U2978 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_45_), 
        .B0(n232), .B1(Input2[45]), .Y(n2915) );
  CLKINVX1 U2979 ( .A(n900), .Y(n899) );
  OAI2B2X1 U2980 ( .A1N(Output2[45]), .A0(n2894), .B0(n2916), .B1(n2895), .Y(
        n900) );
  CLKINVX1 U2981 ( .A(Input2[45]), .Y(n2916) );
  XOR2X1 U2982 ( .A(n2917), .B(n1205), .Y(Output2[45]) );
  CLKINVX1 U2983 ( .A(n2918), .Y(n1205) );
  OAI221X1 U2984 ( .A0(n2919), .A1(n2273), .B0(n2730), .B1(n2229), .C0(n2920), 
        .Y(n2918) );
  MXI2X1 U2985 ( .A(n2921), .B(n2922), .S0(n2923), .Y(n2920) );
  NOR2X1 U2986 ( .A(n2230), .B(n2107), .Y(n2923) );
  OAI22X1 U2987 ( .A0(n2722), .A1(n2645), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[40]), .B1(n2255), .Y(n2922) );
  OAI2BB2X1 U2988 ( .B0(n2255), .B1(n2924), .A0N(n2645), .A1N(n2258), .Y(n2921) );
  XNOR2X1 U2989 ( .A(n2925), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[88]), .Y(
        n2645) );
  XOR2X1 U2990 ( .A(n2926), .B(n2927), .Y(n2919) );
  XOR2X1 U2991 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[80]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[56]), .Y(n2927) );
  CLKNAND2X2 U2992 ( .A(Input2[45]), .B(n2288), .Y(n2917) );
  OAI221X1 U2993 ( .A0(n903), .A1(n178), .B0(n2928), .B1(n149), .C0(n2929), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_44_N3) );
  AOI22XL U2994 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_44_), 
        .B0(n232), .B1(Input2[44]), .Y(n2929) );
  CLKINVX1 U2995 ( .A(n1207), .Y(n2928) );
  CLKINVX1 U2996 ( .A(n904), .Y(n903) );
  OAI2B2X1 U2997 ( .A1N(Output2[44]), .A0(n2894), .B0(n2930), .B1(n2895), .Y(
        n904) );
  XOR2X1 U2998 ( .A(n1207), .B(n2931), .Y(Output2[44]) );
  NOR2X1 U2999 ( .A(n247), .B(n2930), .Y(n2931) );
  CLKINVX1 U3000 ( .A(Input2[44]), .Y(n2930) );
  OAI221X1 U3001 ( .A0(n2230), .A1(n2274), .B0(n276), .B1(n2106), .C0(n2932), 
        .Y(n1207) );
  AOI22XL U3002 ( .A0(n263), .A1(n2933), .B0(n295), .B1(n2934), .Y(n2932) );
  XOR2X1 U3003 ( .A(n2786), .B(n2935), .Y(n2933) );
  XOR2X1 U3004 ( .A(n2430), .B(n2195), .Y(n2935) );
  XNOR2X1 U3005 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_21_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[83]), .Y(n2195) );
  CLKINVX1 U3006 ( .A(n2218), .Y(n2786) );
  MXI2X1 U3007 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[43]), .B(n2656), .S0(
        n308), .Y(n2230) );
  XOR2X1 U3008 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[27]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[91]), .Y(n2656) );
  OAI221X1 U3009 ( .A0(n907), .A1(n178), .B0(n2936), .B1(n149), .C0(n2937), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_43_N3) );
  AOI22XL U3010 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_43_), 
        .B0(n232), .B1(Input2[43]), .Y(n2937) );
  CLKINVX1 U3011 ( .A(n1209), .Y(n2936) );
  CLKINVX1 U3012 ( .A(n908), .Y(n907) );
  OAI2B2X1 U3013 ( .A1N(Output2[43]), .A0(n2894), .B0(n2938), .B1(n2895), .Y(
        n908) );
  XOR2X1 U3014 ( .A(n1209), .B(n2939), .Y(Output2[43]) );
  NOR2X1 U3015 ( .A(n247), .B(n2938), .Y(n2939) );
  CLKINVX1 U3016 ( .A(Input2[43]), .Y(n2938) );
  OAI211XL U3017 ( .A0(n2666), .A1(n2722), .B0(n2940), .C0(n2941), .Y(n1209)
         );
  AOI22XL U3018 ( .A0(n263), .A1(n2942), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[42]), .B1(n2312), .Y(n2941) );
  XOR2X1 U3019 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_11_), .B(n2943), 
        .Y(n2942) );
  XOR2X1 U3020 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[57]), .Y(n2943) );
  MXI2X1 U3021 ( .A(n2944), .B(n2945), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[44]), .Y(n2940) );
  OAI21X1 U3022 ( .A0(n2946), .A1(n279), .B0(n2267), .Y(n2945) );
  NOR2X1 U3023 ( .A(n2106), .B(n2229), .Y(n2946) );
  NOR3X1 U3024 ( .A(n2229), .B(n276), .C(n2106), .Y(n2944) );
  XNOR2X1 U3025 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[26]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[90]), .Y(n2666) );
  OAI221X1 U3026 ( .A0(n911), .A1(n178), .B0(n2947), .B1(n149), .C0(n2948), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_42_N3) );
  AOI22XL U3027 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_42_), 
        .B0(n232), .B1(Input2[42]), .Y(n2948) );
  CLKINVX1 U3028 ( .A(n1211), .Y(n2947) );
  CLKINVX1 U3029 ( .A(n912), .Y(n911) );
  OAI2B2X1 U3030 ( .A1N(Output2[42]), .A0(n2894), .B0(n2949), .B1(n2895), .Y(
        n912) );
  XOR2X1 U3031 ( .A(n1211), .B(n2950), .Y(Output2[42]) );
  NOR2X1 U3032 ( .A(n247), .B(n2949), .Y(n2950) );
  CLKINVX1 U3033 ( .A(Input2[42]), .Y(n2949) );
  OAI221X1 U3034 ( .A0(n2951), .A1(n2273), .B0(n2104), .B1(n2274), .C0(n2952), 
        .Y(n1211) );
  MXI2X1 U3035 ( .A(n2953), .B(n2954), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[40]), .Y(n2952) );
  OAI21X1 U3036 ( .A0(n2955), .A1(n279), .B0(n2267), .Y(n2954) );
  NOR2X1 U3037 ( .A(n2232), .B(n2109), .Y(n2955) );
  NOR3X1 U3038 ( .A(n274), .B(n2232), .C(n2109), .Y(n2953) );
  MXI2X1 U3039 ( .A(n2934), .B(n2681), .S0(n308), .Y(n2104) );
  XOR2X1 U3040 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[92]), .Y(n2681) );
  XNOR2X1 U3041 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_11_), .B(n2106), .Y(
        n2934) );
  XOR2X1 U3042 ( .A(n2956), .B(n2957), .Y(n2951) );
  XOR2X1 U3043 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[84]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[42]), .Y(n2957) );
  OAI221X1 U3044 ( .A0(n915), .A1(n178), .B0(n1212), .B1(n152), .C0(n2958), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_41_N3) );
  AOI22XL U3045 ( .A0(n204), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_41_), 
        .B0(n231), .B1(Input2[41]), .Y(n2958) );
  CLKINVX1 U3046 ( .A(n916), .Y(n915) );
  OAI2B2X1 U3047 ( .A1N(Output2[41]), .A0(n2894), .B0(n2959), .B1(n2895), .Y(
        n916) );
  CLKINVX1 U3048 ( .A(Input2[41]), .Y(n2959) );
  XOR2X1 U3049 ( .A(n2960), .B(n1212), .Y(Output2[41]) );
  CLKINVX1 U3050 ( .A(n2961), .Y(n1212) );
  OAI221X1 U3051 ( .A0(n2962), .A1(n2273), .B0(n2227), .B1(n2274), .C0(n2963), 
        .Y(n2961) );
  AOI22XL U3052 ( .A0(n291), .A1(n2745), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[43]), .B1(n299), .Y(n2963) );
  CLKINVX1 U3053 ( .A(n2232), .Y(n2745) );
  MXI2X1 U3054 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[47]), .B(n2690), .S0(
        n309), .Y(n2227) );
  XOR2X1 U3055 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[31]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[95]), .Y(n2690) );
  XOR2X1 U3056 ( .A(n2964), .B(n2965), .Y(n2962) );
  XOR2X1 U3057 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[87]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[63]), .Y(n2965) );
  CLKNAND2X2 U3058 ( .A(Input2[41]), .B(n2288), .Y(n2960) );
  OAI221X1 U3059 ( .A0(n919), .A1(n177), .B0(n2966), .B1(n149), .C0(n2967), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_40_N3) );
  AOI22XL U3060 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_40_), 
        .B0(n231), .B1(Input2[40]), .Y(n2967) );
  CLKINVX1 U3061 ( .A(n1214), .Y(n2966) );
  CLKINVX1 U3062 ( .A(n920), .Y(n919) );
  OAI2B2X1 U3063 ( .A1N(Output2[40]), .A0(n2894), .B0(n2968), .B1(n2895), .Y(
        n920) );
  XOR2X1 U3064 ( .A(n1214), .B(n2969), .Y(Output2[40]) );
  NOR2X1 U3065 ( .A(n247), .B(n2968), .Y(n2969) );
  CLKINVX1 U3066 ( .A(Input2[40]), .Y(n2968) );
  OAI221X1 U3067 ( .A0(n2107), .A1(n2274), .B0(n282), .B1(n2970), .C0(n2971), 
        .Y(n1214) );
  AOI22XL U3068 ( .A0(n263), .A1(n2972), .B0(n294), .B1(n2900), .Y(n2971) );
  XNOR2X1 U3069 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_10_), .B(n2970), .Y(
        n2900) );
  XOR2X1 U3070 ( .A(n2413), .B(n2973), .Y(n2972) );
  XOR2X1 U3071 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_8_), .B(n2974), 
        .Y(n2973) );
  CLKINVX1 U3072 ( .A(n2074), .Y(n2413) );
  XNOR2X1 U3073 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_20_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[82]), .Y(n2074) );
  CLKINVX1 U3074 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[63]), .Y(n2970) );
  MXI2X1 U3075 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[41]), .B(n2698), .S0(
        n309), .Y(n2107) );
  XOR2X1 U3076 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .Y(n2698) );
  OAI221X1 U3077 ( .A0(n1056), .A1(n177), .B0(n1277), .B1(n149), .C0(n2975), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_4_N3) );
  AOI22XL U3078 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_4_), 
        .B0(n231), .B1(Input2[4]), .Y(n2975) );
  AOI22XL U3079 ( .A0(Input2[4]), .A1(n2627), .B0(n1989), .B1(Output2[4]), .Y(
        n1056) );
  XOR2X1 U3080 ( .A(n2976), .B(n1277), .Y(Output2[4]) );
  AOI221XL U3081 ( .A0(n2977), .A1(n296), .B0(n2873), .B1(n2293), .C0(n2978), 
        .Y(n1277) );
  OAI2BB2X1 U3082 ( .B0(n2024), .B1(n284), .A0N(n2979), .A1N(n269), .Y(n2978)
         );
  CLKINVX1 U3083 ( .A(n2165), .Y(n2873) );
  MXI2X1 U3084 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[3]), .B(n2980), .S0(
        n309), .Y(n2165) );
  XOR2X1 U3085 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[11]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[107]), .Y(n2980) );
  CLKNAND2X2 U3086 ( .A(Input2[4]), .B(n2288), .Y(n2976) );
  OAI221X1 U3087 ( .A0(n2981), .A1(n2300), .B0(n2982), .B1(n2302), .C0(n2983), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_39_N3) );
  AOI22XL U3088 ( .A0(n186), .A1(n923), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1216), .Y(n2983) );
  OAI2B2X1 U3089 ( .A1N(Output2[39]), .A0(n2984), .B0(n2982), .B1(n2985), .Y(
        n923) );
  XOR2X1 U3090 ( .A(n1216), .B(n2986), .Y(Output2[39]) );
  NOR2X1 U3091 ( .A(n247), .B(n2982), .Y(n2986) );
  OAI221X1 U3092 ( .A0(n2116), .A1(n277), .B0(n2267), .B1(n2987), .C0(n2988), 
        .Y(n1216) );
  AOI222XL U3093 ( .A0(n2258), .A1(n2314), .B0(n260), .B1(n2989), .C0(n2312), 
        .C1(n2990), .Y(n2988) );
  XOR2X1 U3094 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_31_), .B(n2991), 
        .Y(n2989) );
  XOR2X1 U3095 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[72]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[39]), .Y(n2991) );
  XOR2X1 U3096 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[80]), .Y(n2314) );
  CLKINVX1 U3097 ( .A(Input2[39]), .Y(n2982) );
  CLKINVX1 U3098 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_39_), .Y(n2981) );
  OAI221X1 U3099 ( .A0(n926), .A1(n177), .B0(n1217), .B1(n149), .C0(n2992), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_38_N3) );
  AOI22XL U3100 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_38_), 
        .B0(n231), .B1(Input2[38]), .Y(n2992) );
  CLKINVX1 U3101 ( .A(n927), .Y(n926) );
  OAI2B2X1 U3102 ( .A1N(Output2[38]), .A0(n2984), .B0(n2993), .B1(n2985), .Y(
        n927) );
  CLKINVX1 U3103 ( .A(Input2[38]), .Y(n2993) );
  XOR2X1 U3104 ( .A(n2994), .B(n1217), .Y(Output2[38]) );
  CLKINVX1 U3105 ( .A(n2995), .Y(n1217) );
  OAI211XL U3106 ( .A0(n285), .A1(n2987), .B0(n2996), .C0(n2997), .Y(n2995) );
  AOI22XL U3107 ( .A0(n263), .A1(n2998), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[34]), .B1(n299), .Y(n2997) );
  XOR2X1 U3108 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_), .B(n2999), 
        .Y(n2998) );
  XOR2X1 U3109 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[76]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .Y(n2999) );
  MXI2X1 U3110 ( .A(n3000), .B(n3001), .S0(n3002), .Y(n2996) );
  NOR2X1 U3111 ( .A(n2111), .B(n2234), .Y(n3002) );
  OAI22X1 U3112 ( .A0(n2722), .A1(n2327), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[36]), .B1(n2255), .Y(n3001) );
  OAI2BB2X1 U3113 ( .B0(n2255), .B1(n3003), .A0N(n2327), .A1N(n2258), .Y(n3000) );
  XNOR2X1 U3114 ( .A(n3004), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[84]), .Y(
        n2327) );
  CLKNAND2X2 U3115 ( .A(Input2[38]), .B(n2288), .Y(n2994) );
  OAI221X1 U3116 ( .A0(n930), .A1(n177), .B0(n1218), .B1(n149), .C0(n3005), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_37_N3) );
  AOI22XL U3117 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_37_), 
        .B0(n231), .B1(Input2[37]), .Y(n3005) );
  CLKINVX1 U3118 ( .A(n931), .Y(n930) );
  OAI2B2X1 U3119 ( .A1N(Output2[37]), .A0(n2984), .B0(n3006), .B1(n2985), .Y(
        n931) );
  CLKINVX1 U3120 ( .A(Input2[37]), .Y(n3006) );
  XOR2X1 U3121 ( .A(n3007), .B(n1218), .Y(Output2[37]) );
  CLKINVX1 U3122 ( .A(n3008), .Y(n1218) );
  OAI221X1 U3123 ( .A0(n3009), .A1(n2273), .B0(n2730), .B1(n2236), .C0(n3010), 
        .Y(n3008) );
  MXI2X1 U3124 ( .A(n3011), .B(n3012), .S0(n3013), .Y(n3010) );
  NOR2X1 U3125 ( .A(n2237), .B(n2114), .Y(n3013) );
  OAI22X1 U3126 ( .A0(n2722), .A1(n2340), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[32]), .B1(n2255), .Y(n3012) );
  OAI2BB2X1 U3127 ( .B0(n2255), .B1(n3014), .A0N(n2340), .A1N(n2258), .Y(n3011) );
  XNOR2X1 U3128 ( .A(n3015), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[80]), .Y(
        n2340) );
  XOR2X1 U3129 ( .A(n3016), .B(n3017), .Y(n3009) );
  XOR2X1 U3130 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[72]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .Y(n3017) );
  CLKNAND2X2 U3131 ( .A(Input2[37]), .B(n2288), .Y(n3007) );
  OAI221X1 U3132 ( .A0(n934), .A1(n177), .B0(n3018), .B1(n148), .C0(n3019), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_36_N3) );
  AOI22XL U3133 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_36_), 
        .B0(n231), .B1(Input2[36]), .Y(n3019) );
  CLKINVX1 U3134 ( .A(n1220), .Y(n3018) );
  CLKINVX1 U3135 ( .A(n935), .Y(n934) );
  OAI2B2X1 U3136 ( .A1N(Output2[36]), .A0(n2984), .B0(n3020), .B1(n2985), .Y(
        n935) );
  XOR2X1 U3137 ( .A(n1220), .B(n3021), .Y(Output2[36]) );
  NOR2X1 U3138 ( .A(n247), .B(n3020), .Y(n3021) );
  CLKINVX1 U3139 ( .A(Input2[36]), .Y(n3020) );
  OAI221X1 U3140 ( .A0(n2237), .A1(n2274), .B0(n284), .B1(n2113), .C0(n3022), 
        .Y(n1220) );
  AOI22XL U3141 ( .A0(n264), .A1(n3023), .B0(n295), .B1(n3024), .Y(n3022) );
  XNOR2X1 U3142 ( .A(n2225), .B(n3025), .Y(n3023) );
  XOR2X1 U3143 ( .A(n2531), .B(n2203), .Y(n3025) );
  XNOR2X1 U3144 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_19_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[75]), .Y(n2203) );
  MXI2X1 U3145 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[35]), .B(n2351), .S0(
        n309), .Y(n2237) );
  XOR2X1 U3146 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[19]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[83]), .Y(n2351) );
  OAI221X1 U3147 ( .A0(n938), .A1(n177), .B0(n3026), .B1(n148), .C0(n3027), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_35_N3) );
  AOI22XL U3148 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_35_), 
        .B0(n231), .B1(Input2[35]), .Y(n3027) );
  CLKINVX1 U3149 ( .A(n1222), .Y(n3026) );
  CLKINVX1 U3150 ( .A(n939), .Y(n938) );
  OAI2B2X1 U3151 ( .A1N(Output2[35]), .A0(n2984), .B0(n3028), .B1(n2985), .Y(
        n939) );
  XOR2X1 U3152 ( .A(n1222), .B(n3029), .Y(Output2[35]) );
  NOR2X1 U3153 ( .A(n247), .B(n3028), .Y(n3029) );
  CLKINVX1 U3154 ( .A(Input2[35]), .Y(n3028) );
  OAI211XL U3155 ( .A0(n2361), .A1(n2722), .B0(n3030), .C0(n3031), .Y(n1222)
         );
  AOI22XL U3156 ( .A0(n262), .A1(n3032), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[34]), .B1(n2312), .Y(n3031) );
  XOR2X1 U3157 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_27_), .B(n3033), 
        .Y(n3032) );
  XOR2X1 U3158 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[73]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[49]), .Y(n3033) );
  MXI2X1 U3159 ( .A(n3034), .B(n3035), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[36]), .Y(n3030) );
  OAI21X1 U3160 ( .A0(n3036), .A1(n279), .B0(n2267), .Y(n3035) );
  NOR2X1 U3161 ( .A(n2113), .B(n2236), .Y(n3036) );
  NOR3X1 U3162 ( .A(n2236), .B(n276), .C(n2113), .Y(n3034) );
  XNOR2X1 U3163 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[18]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[82]), .Y(n2361) );
  OAI221X1 U3164 ( .A0(n942), .A1(n177), .B0(n3037), .B1(n148), .C0(n3038), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_34_N3) );
  AOI22XL U3165 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_34_), 
        .B0(n231), .B1(Input2[34]), .Y(n3038) );
  CLKINVX1 U3166 ( .A(n1224), .Y(n3037) );
  CLKINVX1 U3167 ( .A(n943), .Y(n942) );
  OAI2B2X1 U3168 ( .A1N(Output2[34]), .A0(n2984), .B0(n3039), .B1(n2985), .Y(
        n943) );
  XOR2X1 U3169 ( .A(n1224), .B(n3040), .Y(Output2[34]) );
  NOR2X1 U3170 ( .A(n247), .B(n3039), .Y(n3040) );
  CLKINVX1 U3171 ( .A(Input2[34]), .Y(n3039) );
  OAI221X1 U3172 ( .A0(n3041), .A1(n2273), .B0(n2111), .B1(n2274), .C0(n3042), 
        .Y(n1224) );
  MXI2X1 U3173 ( .A(n3043), .B(n3044), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[32]), .Y(n3042) );
  OAI21X1 U3174 ( .A0(n3045), .A1(n280), .B0(n2267), .Y(n3044) );
  NOR2X1 U3175 ( .A(n2239), .B(n2116), .Y(n3045) );
  NOR3X1 U3176 ( .A(n274), .B(n2239), .C(n2116), .Y(n3043) );
  MXI2X1 U3177 ( .A(n3024), .B(n2376), .S0(n309), .Y(n2111) );
  XOR2X1 U3178 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[84]), .Y(n2376) );
  XNOR2X1 U3179 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_9_), .B(n2113), .Y(
        n3024) );
  XOR2X1 U3180 ( .A(n3046), .B(n3047), .Y(n3041) );
  XOR2X1 U3181 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[76]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[34]), .Y(n3047) );
  OAI221X1 U3182 ( .A0(n946), .A1(n177), .B0(n1225), .B1(n148), .C0(n3048), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_33_N3) );
  AOI22XL U3183 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_33_), 
        .B0(n231), .B1(Input2[33]), .Y(n3048) );
  CLKINVX1 U3184 ( .A(n947), .Y(n946) );
  OAI2B2X1 U3185 ( .A1N(Output2[33]), .A0(n2984), .B0(n3049), .B1(n2985), .Y(
        n947) );
  CLKINVX1 U3186 ( .A(Input2[33]), .Y(n3049) );
  XOR2X1 U3187 ( .A(n3050), .B(n1225), .Y(Output2[33]) );
  CLKINVX1 U3188 ( .A(n3051), .Y(n1225) );
  OAI221X1 U3189 ( .A0(n3052), .A1(n2273), .B0(n2234), .B1(n2274), .C0(n3053), 
        .Y(n3051) );
  AOI22XL U3190 ( .A0(n291), .A1(n2839), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[35]), .B1(n300), .Y(n3053) );
  CLKINVX1 U3191 ( .A(n2239), .Y(n2839) );
  MXI2X1 U3192 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[39]), .B(n2394), .S0(
        n309), .Y(n2234) );
  XOR2X1 U3193 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[23]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[87]), .Y(n2394) );
  XOR2X1 U3194 ( .A(n3054), .B(n3055), .Y(n3052) );
  XOR2X1 U3195 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[79]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[55]), .Y(n3055) );
  CLKNAND2X2 U3196 ( .A(Input2[33]), .B(n2288), .Y(n3050) );
  OAI221X1 U3197 ( .A0(n950), .A1(n177), .B0(n3056), .B1(n148), .C0(n3057), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_32_N3) );
  AOI22XL U3198 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_32_), 
        .B0(n231), .B1(Input2[32]), .Y(n3057) );
  CLKINVX1 U3199 ( .A(n1227), .Y(n3056) );
  CLKINVX1 U3200 ( .A(n951), .Y(n950) );
  OAI2B2X1 U3201 ( .A1N(Output2[32]), .A0(n2984), .B0(n3058), .B1(n2985), .Y(
        n951) );
  XOR2X1 U3202 ( .A(n1227), .B(n3059), .Y(Output2[32]) );
  NOR2X1 U3203 ( .A(n247), .B(n3058), .Y(n3059) );
  CLKINVX1 U3204 ( .A(Input2[32]), .Y(n3058) );
  OAI221X1 U3205 ( .A0(n2114), .A1(n2274), .B0(n276), .B1(n3060), .C0(n3061), 
        .Y(n1227) );
  AOI22XL U3206 ( .A0(n264), .A1(n3062), .B0(n295), .B1(n2990), .Y(n3061) );
  XNOR2X1 U3207 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_8_), .B(n3060), .Y(
        n2990) );
  XOR2X1 U3208 ( .A(n2513), .B(n3063), .Y(n3062) );
  XOR2X1 U3209 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_24_), .B(n3064), 
        .Y(n3063) );
  CLKINVX1 U3210 ( .A(n2081), .Y(n2513) );
  XNOR2X1 U3211 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_18_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[74]), .Y(n2081) );
  MXI2X1 U3212 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[33]), .B(n2402), .S0(
        n309), .Y(n2114) );
  XOR2X1 U3213 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .Y(n2402) );
  OAI221X1 U3214 ( .A0(n3065), .A1(n2300), .B0(n3066), .B1(n2302), .C0(n3067), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_31_N3) );
  AOI22XL U3215 ( .A0(n186), .A1(n954), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1229), .Y(n3067) );
  OAI2B2X1 U3216 ( .A1N(Output2[31]), .A0(n3068), .B0(n3066), .B1(n3069), .Y(
        n954) );
  XOR2X1 U3217 ( .A(n1229), .B(n3070), .Y(Output2[31]) );
  NOR2X1 U3218 ( .A(n247), .B(n3066), .Y(n3070) );
  OAI221X1 U3219 ( .A0(n3071), .A1(n2273), .B0(n2267), .B1(n3072), .C0(n3073), 
        .Y(n1229) );
  AOI222XL U3220 ( .A0(n291), .A1(n2298), .B0(n2258), .B1(n3074), .C0(n2312), 
        .C1(n3075), .Y(n3073) );
  XOR2X1 U3221 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[96]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]), .Y(n3074) );
  CLKINVX1 U3222 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .Y(n3072) );
  CLKINVX1 U3223 ( .A(Input2[31]), .Y(n3066) );
  CLKINVX1 U3224 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_31_), .Y(n3065) );
  OAI221X1 U3225 ( .A0(n957), .A1(n177), .B0(n1230), .B1(n148), .C0(n3076), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_30_N3) );
  AOI22XL U3226 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_30_), 
        .B0(n231), .B1(Input2[30]), .Y(n3076) );
  CLKINVX1 U3227 ( .A(n958), .Y(n957) );
  OAI2B2X1 U3228 ( .A1N(Output2[30]), .A0(n3068), .B0(n3077), .B1(n3069), .Y(
        n958) );
  CLKINVX1 U3229 ( .A(Input2[30]), .Y(n3077) );
  XOR2X1 U3230 ( .A(n3078), .B(n1230), .Y(Output2[30]) );
  CLKINVX1 U3231 ( .A(n3079), .Y(n1230) );
  OAI221X1 U3232 ( .A0(n3080), .A1(n2274), .B0(n3081), .B1(n2273), .C0(n3082), 
        .Y(n3079) );
  AOI22XL U3233 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[26]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .B1(n292), .Y(n3082) );
  XOR2X1 U3234 ( .A(n3083), .B(n3084), .Y(n3080) );
  MXI2X1 U3235 ( .A(n2914), .B(n3085), .S0(n309), .Y(n3084) );
  XOR2X1 U3236 ( .A(n3086), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[4]), .Y(
        n3085) );
  CLKINVX1 U3237 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[28]), .Y(n2914) );
  OR2X1 U3238 ( .A(n2241), .B(n2118), .Y(n3083) );
  CLKNAND2X2 U3239 ( .A(Input2[30]), .B(n2288), .Y(n3078) );
  OAI221X1 U3240 ( .A0(n1059), .A1(n177), .B0(n3087), .B1(n148), .C0(n3088), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_3_N3) );
  AOI22XL U3241 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_3_), 
        .B0(n231), .B1(Input2[3]), .Y(n3088) );
  CLKINVX1 U3242 ( .A(n1279), .Y(n3087) );
  AOI22XL U3243 ( .A0(n1989), .A1(Output2[3]), .B0(Input2[3]), .B1(n2627), .Y(
        n1059) );
  XOR2X1 U3244 ( .A(n1279), .B(n3089), .Y(Output2[3]) );
  NOR2BX1 U3245 ( .AN(Input2[3]), .B(n254), .Y(n3089) );
  OAI2B11X1 U3246 ( .A1N(n2262), .A0(n2273), .B0(n3090), .C0(n3091), .Y(n1279)
         );
  AOI22XL U3247 ( .A0(n2258), .A1(n3092), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[2]), .B1(n2312), .Y(n3091) );
  XOR2X1 U3248 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[106]), .Y(n3092) );
  MXI2X1 U3249 ( .A(n3093), .B(n3094), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[4]), .Y(n3090) );
  OAI21X1 U3250 ( .A0(n3095), .A1(n280), .B0(n2267), .Y(n3094) );
  NOR2X1 U3251 ( .A(n2024), .B(n2143), .Y(n3095) );
  NOR3X1 U3252 ( .A(n2143), .B(n276), .C(n2024), .Y(n3093) );
  CLKINVX1 U3253 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]), .Y(n2024) );
  CLKINVX1 U3254 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[7]), .Y(n2143) );
  XOR2X1 U3255 ( .A(n2804), .B(n2662), .Y(n2262) );
  XOR2X1 U3256 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_19_), .B(n3096), 
        .Y(n2662) );
  CLKINVX1 U3257 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[49]), .Y(n2804) );
  OAI221X1 U3258 ( .A0(n961), .A1(n177), .B0(n3097), .B1(n148), .C0(n3098), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_29_N3) );
  AOI22XL U3259 ( .A0(n203), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_29_), 
        .B0(n231), .B1(Input2[29]), .Y(n3098) );
  CLKINVX1 U3260 ( .A(n1232), .Y(n3097) );
  CLKINVX1 U3261 ( .A(n962), .Y(n961) );
  OAI2B2X1 U3262 ( .A1N(Output2[29]), .A0(n3068), .B0(n3099), .B1(n3069), .Y(
        n962) );
  XOR2X1 U3263 ( .A(n1232), .B(n3100), .Y(Output2[29]) );
  NOR2X1 U3264 ( .A(n248), .B(n3099), .Y(n3100) );
  CLKINVX1 U3265 ( .A(Input2[29]), .Y(n3099) );
  OAI222X1 U3266 ( .A0(n2730), .A1(n2243), .B0(n3101), .B1(n2274), .C0(n3102), 
        .C1(n2273), .Y(n1232) );
  XOR2X1 U3267 ( .A(n3103), .B(n3104), .Y(n3101) );
  MXI2X1 U3268 ( .A(n2925), .B(n3105), .S0(n309), .Y(n3104) );
  XOR2X1 U3269 ( .A(n2829), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[96]), .Y(
        n3105) );
  CLKINVX1 U3270 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[0]), .Y(n2829) );
  CLKINVX1 U3271 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[24]), .Y(n2925) );
  CLKNAND2X2 U3272 ( .A(n3106), .B(n3107), .Y(n3103) );
  OAI221X1 U3273 ( .A0(n965), .A1(n176), .B0(n1234), .B1(n148), .C0(n3108), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_28_N3) );
  AOI22XL U3274 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_28_), 
        .B0(n230), .B1(Input2[28]), .Y(n3108) );
  CLKINVX1 U3275 ( .A(n966), .Y(n965) );
  OAI2B2X1 U3276 ( .A1N(Input2[28]), .A0(n3069), .B0(n3109), .B1(n3068), .Y(
        n966) );
  CLKINVX1 U3277 ( .A(Output2[28]), .Y(n3109) );
  XOR2X1 U3278 ( .A(n3110), .B(n1234), .Y(Output2[28]) );
  AOI221XL U3279 ( .A0(n3111), .A1(n296), .B0(n3107), .B1(n2293), .C0(n3112), 
        .Y(n1234) );
  OAI2BB2X1 U3280 ( .B0(n2120), .B1(n284), .A0N(n3113), .A1N(n268), .Y(n3112)
         );
  CLKINVX1 U3281 ( .A(n2121), .Y(n3107) );
  MXI2X1 U3282 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[27]), .B(n3114), .S0(
        n309), .Y(n2121) );
  XOR2X1 U3283 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[99]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[3]), .Y(n3114) );
  CLKNAND2X2 U3284 ( .A(Input2[28]), .B(n2288), .Y(n3110) );
  OAI221X1 U3285 ( .A0(n969), .A1(n176), .B0(n3115), .B1(n148), .C0(n3116), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_27_N3) );
  AOI22XL U3286 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_27_), 
        .B0(n230), .B1(Input2[27]), .Y(n3116) );
  CLKINVX1 U3287 ( .A(n1236), .Y(n3115) );
  CLKINVX1 U3288 ( .A(n970), .Y(n969) );
  OAI2B2X1 U3289 ( .A1N(Output2[27]), .A0(n3068), .B0(n3117), .B1(n3069), .Y(
        n970) );
  XOR2X1 U3290 ( .A(n1236), .B(n3118), .Y(Output2[27]) );
  NOR2X1 U3291 ( .A(n248), .B(n3117), .Y(n3118) );
  CLKINVX1 U3292 ( .A(Input2[27]), .Y(n3117) );
  OAI2B11X1 U3293 ( .A1N(n3119), .A0(n2273), .B0(n3120), .C0(n3121), .Y(n1236)
         );
  AOI22XL U3294 ( .A0(n2258), .A1(n3122), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[26]), .B1(n2312), .Y(n3121) );
  XOR2X1 U3295 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[98]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[2]), .Y(n3122) );
  MXI2X1 U3296 ( .A(n3123), .B(n3124), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[28]), .Y(n3120) );
  OAI21X1 U3297 ( .A0(n3125), .A1(n280), .B0(n2267), .Y(n3124) );
  NOR2X1 U3298 ( .A(n2120), .B(n2243), .Y(n3125) );
  NOR3X1 U3299 ( .A(n2243), .B(n276), .C(n2120), .Y(n3123) );
  CLKINVX1 U3300 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]), .Y(n2120) );
  CLKINVX1 U3301 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[31]), .Y(n2243) );
  OAI221X1 U3302 ( .A0(n973), .A1(n176), .B0(n3126), .B1(n148), .C0(n3127), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_26_N3) );
  AOI22XL U3303 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_26_), 
        .B0(n230), .B1(Input2[26]), .Y(n3127) );
  CLKINVX1 U3304 ( .A(n1238), .Y(n3126) );
  CLKINVX1 U3305 ( .A(n974), .Y(n973) );
  OAI2B2X1 U3306 ( .A1N(Output2[26]), .A0(n3068), .B0(n3128), .B1(n3069), .Y(
        n974) );
  XOR2X1 U3307 ( .A(n1238), .B(n3129), .Y(Output2[26]) );
  NOR2X1 U3308 ( .A(n248), .B(n3128), .Y(n3129) );
  CLKINVX1 U3309 ( .A(Input2[26]), .Y(n3128) );
  OAI221X1 U3310 ( .A0(n2118), .A1(n2274), .B0(n3130), .B1(n2273), .C0(n3131), 
        .Y(n1238) );
  MXI2X1 U3311 ( .A(n3132), .B(n3133), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[24]), .Y(n3131) );
  OAI21X1 U3312 ( .A0(n3134), .A1(n280), .B0(n2267), .Y(n3133) );
  NOR2X1 U3313 ( .A(n2006), .B(n2123), .Y(n3134) );
  NOR3X1 U3314 ( .A(n274), .B(n2006), .C(n2123), .Y(n3132) );
  CLKINVX1 U3315 ( .A(n2298), .Y(n2006) );
  XOR2X1 U3316 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_6_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[26]), .Y(n2298) );
  MXI2X1 U3317 ( .A(n3111), .B(n3135), .S0(n309), .Y(n2118) );
  XOR2X1 U3318 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[100]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]), .Y(n3135) );
  XOR2X1 U3319 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_7_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]), .Y(n3111) );
  OAI221X1 U3320 ( .A0(n977), .A1(n176), .B0(n1239), .B1(n148), .C0(n3136), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_25_N3) );
  AOI22XL U3321 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_25_), 
        .B0(n230), .B1(Input2[25]), .Y(n3136) );
  CLKINVX1 U3322 ( .A(n978), .Y(n977) );
  OAI2B2X1 U3323 ( .A1N(Output2[25]), .A0(n3068), .B0(n3137), .B1(n3069), .Y(
        n978) );
  CLKINVX1 U3324 ( .A(Input2[25]), .Y(n3137) );
  XOR2X1 U3325 ( .A(n3138), .B(n1239), .Y(Output2[25]) );
  CLKINVX1 U3326 ( .A(n3139), .Y(n1239) );
  OAI221X1 U3327 ( .A0(n2241), .A1(n2274), .B0(n3140), .B1(n2273), .C0(n3141), 
        .Y(n3139) );
  AOI2BB2X1 U3328 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[27]), .B1(n294), 
        .A0N(n285), .A1N(n2123), .Y(n3141) );
  MXI2X1 U3329 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[31]), .B(n3142), .S0(
        n309), .Y(n2241) );
  XOR2X1 U3330 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[7]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[103]), .Y(n3142) );
  CLKNAND2X2 U3331 ( .A(Input2[25]), .B(n2288), .Y(n3138) );
  OAI221X1 U3332 ( .A0(n981), .A1(n176), .B0(n1241), .B1(n148), .C0(n3143), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_24_N3) );
  AOI22XL U3333 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_24_), 
        .B0(n230), .B1(Input2[24]), .Y(n3143) );
  CLKINVX1 U3334 ( .A(n982), .Y(n981) );
  OAI2B2X1 U3335 ( .A1N(Input2[24]), .A0(n3069), .B0(n3144), .B1(n3068), .Y(
        n982) );
  CLKINVX1 U3336 ( .A(Output2[24]), .Y(n3144) );
  XOR2X1 U3337 ( .A(n3145), .B(n1241), .Y(Output2[24]) );
  AOI221XL U3338 ( .A0(n3075), .A1(n296), .B0(n3106), .B1(n2293), .C0(n3146), 
        .Y(n1241) );
  AO22X1 U3339 ( .A0(n266), .A1(n3147), .B0(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]), .B1(n292), .Y(n3146) );
  CLKINVX1 U3340 ( .A(n2003), .Y(n3106) );
  MXI2X1 U3341 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .B(n3148), .S0(
        n310), .Y(n2003) );
  XOR2X1 U3342 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[97]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .Y(n3148) );
  XOR2X1 U3343 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_6_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]), .Y(n3075) );
  CLKNAND2X2 U3344 ( .A(Input2[24]), .B(n2288), .Y(n3145) );
  OAI221X1 U3345 ( .A0(n3149), .A1(n2300), .B0(n3150), .B1(n2302), .C0(n3151), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_23_N3) );
  AOI22XL U3346 ( .A0(n186), .A1(n985), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1243), .Y(n3151) );
  OAI2B2X1 U3347 ( .A1N(Output2[23]), .A0(n3152), .B0(n3150), .B1(n3153), .Y(
        n985) );
  XOR2X1 U3348 ( .A(n1243), .B(n3154), .Y(Output2[23]) );
  NOR2X1 U3349 ( .A(n248), .B(n3150), .Y(n3154) );
  OAI221X1 U3350 ( .A0(n3155), .A1(n2273), .B0(n2267), .B1(n3156), .C0(n3157), 
        .Y(n1243) );
  AOI222XL U3351 ( .A0(n291), .A1(n3158), .B0(n2258), .B1(n3159), .C0(n2312), 
        .C1(n3160), .Y(n3157) );
  XOR2X1 U3352 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[120]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]), .Y(n3159) );
  CLKINVX1 U3353 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .Y(n3156) );
  CLKINVX1 U3354 ( .A(Input2[23]), .Y(n3150) );
  CLKINVX1 U3355 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_23_), .Y(n3149) );
  OAI221X1 U3356 ( .A0(n988), .A1(n176), .B0(n1244), .B1(n148), .C0(n3161), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_22_N3) );
  AOI22XL U3357 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_22_), 
        .B0(n230), .B1(Input2[22]), .Y(n3161) );
  CLKINVX1 U3358 ( .A(n989), .Y(n988) );
  OAI2B2X1 U3359 ( .A1N(Output2[22]), .A0(n3152), .B0(n3162), .B1(n3153), .Y(
        n989) );
  CLKINVX1 U3360 ( .A(Input2[22]), .Y(n3162) );
  XOR2X1 U3361 ( .A(n3163), .B(n1244), .Y(Output2[22]) );
  CLKINVX1 U3362 ( .A(n3164), .Y(n1244) );
  OAI221X1 U3363 ( .A0(n3165), .A1(n2274), .B0(n3166), .B1(n2273), .C0(n3167), 
        .Y(n3164) );
  AOI22XL U3364 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[18]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .B1(n292), .Y(n3167) );
  XOR2X1 U3365 ( .A(n3168), .B(n3169), .Y(n3165) );
  MXI2X1 U3366 ( .A(n3004), .B(n3170), .S0(n310), .Y(n3169) );
  XOR2X1 U3367 ( .A(n3171), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[28]), .Y(
        n3170) );
  CLKINVX1 U3368 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[20]), .Y(n3004) );
  OR2X1 U3369 ( .A(n2125), .B(n2008), .Y(n3168) );
  CLKNAND2X2 U3370 ( .A(Input2[22]), .B(n2288), .Y(n3163) );
  OAI221X1 U3371 ( .A0(n992), .A1(n176), .B0(n3172), .B1(n148), .C0(n3173), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_21_N3) );
  AOI22XL U3372 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_21_), 
        .B0(n230), .B1(Input2[21]), .Y(n3173) );
  CLKINVX1 U3373 ( .A(n1246), .Y(n3172) );
  CLKINVX1 U3374 ( .A(n993), .Y(n992) );
  OAI2B2X1 U3375 ( .A1N(Output2[21]), .A0(n3152), .B0(n3174), .B1(n3153), .Y(
        n993) );
  XOR2X1 U3376 ( .A(n1246), .B(n3175), .Y(Output2[21]) );
  NOR2X1 U3377 ( .A(n248), .B(n3174), .Y(n3175) );
  CLKINVX1 U3378 ( .A(Input2[21]), .Y(n3174) );
  OAI222X1 U3379 ( .A0(n2730), .A1(n2127), .B0(n3176), .B1(n2274), .C0(n3177), 
        .C1(n2273), .Y(n1246) );
  XOR2X1 U3380 ( .A(n3178), .B(n3179), .Y(n3176) );
  MXI2X1 U3381 ( .A(n3015), .B(n3180), .S0(n310), .Y(n3179) );
  XOR2X1 U3382 ( .A(n3181), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[24]), .Y(
        n3180) );
  CLKINVX1 U3383 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[16]), .Y(n3015) );
  CLKNAND2X2 U3384 ( .A(n3182), .B(n3183), .Y(n3178) );
  OAI221X1 U3385 ( .A0(n996), .A1(n176), .B0(n1248), .B1(n148), .C0(n3184), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_20_N3) );
  AOI22XL U3386 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_20_), 
        .B0(n230), .B1(Input2[20]), .Y(n3184) );
  CLKINVX1 U3387 ( .A(n997), .Y(n996) );
  OAI2B2X1 U3388 ( .A1N(Input2[20]), .A0(n3153), .B0(n3185), .B1(n3152), .Y(
        n997) );
  CLKINVX1 U3389 ( .A(Output2[20]), .Y(n3185) );
  XOR2X1 U3390 ( .A(n3186), .B(n1248), .Y(Output2[20]) );
  AOI221XL U3391 ( .A0(n3187), .A1(n296), .B0(n3183), .B1(n2293), .C0(n3188), 
        .Y(n1248) );
  OAI2BB2X1 U3392 ( .B0(n2010), .B1(n284), .A0N(n3189), .A1N(n268), .Y(n3188)
         );
  CLKINVX1 U3393 ( .A(n2129), .Y(n3183) );
  MXI2X1 U3394 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[19]), .B(n3190), .S0(
        n310), .Y(n2129) );
  XOR2X1 U3395 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[27]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[123]), .Y(n3190) );
  CLKNAND2X2 U3396 ( .A(Input2[20]), .B(n2288), .Y(n3186) );
  OAI221X1 U3397 ( .A0(n1062), .A1(n176), .B0(n3191), .B1(n147), .C0(n3192), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_2_N3) );
  AOI22XL U3398 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_2_), 
        .B0(n230), .B1(Input2[2]), .Y(n3192) );
  CLKINVX1 U3399 ( .A(n1281), .Y(n3191) );
  AOI22XL U3400 ( .A0(n1989), .A1(Output2[2]), .B0(Input2[2]), .B1(n2627), .Y(
        n1062) );
  XOR2X1 U3401 ( .A(n1281), .B(n3193), .Y(Output2[2]) );
  NOR2BX1 U3402 ( .AN(Input2[2]), .B(n254), .Y(n3193) );
  OAI221X1 U3403 ( .A0(n2022), .A1(n2274), .B0(n2279), .B1(n2273), .C0(n3194), 
        .Y(n1281) );
  MXI2X1 U3404 ( .A(n3195), .B(n3196), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[0]), .Y(n3194) );
  OAI21X1 U3405 ( .A0(n3197), .A1(n280), .B0(n2267), .Y(n3196) );
  NOR2X1 U3406 ( .A(n2048), .B(n2167), .Y(n3197) );
  NOR3X1 U3407 ( .A(n274), .B(n2048), .C(n2167), .Y(n3195) );
  CLKINVX1 U3408 ( .A(n2632), .Y(n2048) );
  XOR2X1 U3409 ( .A(n2099), .B(n2675), .Y(n2279) );
  XNOR2X1 U3410 ( .A(n3198), .B(Inst_forkAE_CipherInst_RF_S_MID_C2[100]), .Y(
        n2675) );
  CLKINVX1 U3411 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[34]), .Y(n2099) );
  MXI2X1 U3412 ( .A(n2977), .B(n3199), .S0(n310), .Y(n2022) );
  XOR2X1 U3413 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[108]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]), .Y(n3199) );
  XOR2X1 U3414 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_1_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]), .Y(n2977) );
  OAI221X1 U3415 ( .A0(n1000), .A1(n176), .B0(n3200), .B1(n147), .C0(n3201), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_19_N3) );
  AOI22XL U3416 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_19_), 
        .B0(n230), .B1(Input2[19]), .Y(n3201) );
  CLKINVX1 U3417 ( .A(n1250), .Y(n3200) );
  CLKINVX1 U3418 ( .A(n1001), .Y(n1000) );
  OAI2B2X1 U3419 ( .A1N(Output2[19]), .A0(n3152), .B0(n3202), .B1(n3153), .Y(
        n1001) );
  XOR2X1 U3420 ( .A(n1250), .B(n3203), .Y(Output2[19]) );
  NOR2X1 U3421 ( .A(n248), .B(n3202), .Y(n3203) );
  CLKINVX1 U3422 ( .A(Input2[19]), .Y(n3202) );
  OAI2B11X1 U3423 ( .A1N(n3204), .A0(n2273), .B0(n3205), .C0(n3206), .Y(n1250)
         );
  AOI22XL U3424 ( .A0(n2258), .A1(n3207), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[18]), .B1(n2312), .Y(n3206) );
  XOR2X1 U3425 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[26]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[122]), .Y(n3207) );
  MXI2X1 U3426 ( .A(n3208), .B(n3209), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[20]), .Y(n3205) );
  OAI21X1 U3427 ( .A0(n3210), .A1(n281), .B0(n2267), .Y(n3209) );
  NOR2X1 U3428 ( .A(n2127), .B(n2010), .Y(n3210) );
  NOR3X1 U3429 ( .A(n2010), .B(n2127), .C(n278), .Y(n3208) );
  CLKINVX1 U3430 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[23]), .Y(n2127) );
  CLKINVX1 U3431 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]), .Y(n2010) );
  OAI221X1 U3432 ( .A0(n1004), .A1(n176), .B0(n3211), .B1(n147), .C0(n3212), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_18_N3) );
  AOI22XL U3433 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_18_), 
        .B0(n230), .B1(Input2[18]), .Y(n3212) );
  CLKINVX1 U3434 ( .A(n1252), .Y(n3211) );
  CLKINVX1 U3435 ( .A(n1005), .Y(n1004) );
  OAI2B2X1 U3436 ( .A1N(Output2[18]), .A0(n3152), .B0(n3213), .B1(n3153), .Y(
        n1005) );
  XOR2X1 U3437 ( .A(n1252), .B(n3214), .Y(Output2[18]) );
  NOR2X1 U3438 ( .A(n248), .B(n3213), .Y(n3214) );
  CLKINVX1 U3439 ( .A(Input2[18]), .Y(n3213) );
  OAI221X1 U3440 ( .A0(n2008), .A1(n2274), .B0(n3215), .B1(n2273), .C0(n3216), 
        .Y(n1252) );
  MXI2X1 U3441 ( .A(n3217), .B(n3218), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[16]), .Y(n3216) );
  OAI21X1 U3442 ( .A0(n3219), .A1(n280), .B0(n2267), .Y(n3218) );
  NOR2X1 U3443 ( .A(n2013), .B(n2131), .Y(n3219) );
  NOR3X1 U3444 ( .A(n274), .B(n2013), .C(n2131), .Y(n3217) );
  MXI2X1 U3445 ( .A(n3187), .B(n3220), .S0(n310), .Y(n2008) );
  XOR2X1 U3446 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[124]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[2]), .Y(n3220) );
  XOR2X1 U3447 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_5_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]), .Y(n3187) );
  OAI221X1 U3448 ( .A0(n1008), .A1(n176), .B0(n3221), .B1(n147), .C0(n3222), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_17_N3) );
  AOI22XL U3449 ( .A0(n202), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_17_), 
        .B0(n230), .B1(Input2[17]), .Y(n3222) );
  CLKINVX1 U3450 ( .A(n1254), .Y(n3221) );
  CLKINVX1 U3451 ( .A(n1009), .Y(n1008) );
  OAI2B2X1 U3452 ( .A1N(Output2[17]), .A0(n3152), .B0(n3223), .B1(n3153), .Y(
        n1009) );
  XOR2X1 U3453 ( .A(n1254), .B(n3224), .Y(Output2[17]) );
  NOR2X1 U3454 ( .A(n248), .B(n3223), .Y(n3224) );
  CLKINVX1 U3455 ( .A(Input2[17]), .Y(n3223) );
  OAI221X1 U3456 ( .A0(n2125), .A1(n2274), .B0(n2131), .B1(n278), .C0(n3225), 
        .Y(n1254) );
  AOI22XL U3457 ( .A0(n264), .A1(n3226), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[19]), .B1(n299), .Y(n3225) );
  MXI2X1 U3458 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[23]), .B(n3227), .S0(
        n310), .Y(n2125) );
  XOR2X1 U3459 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[31]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[127]), .Y(n3227) );
  OAI221X1 U3460 ( .A0(n1012), .A1(n175), .B0(n1256), .B1(n147), .C0(n3228), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_16_N3) );
  AOI22XL U3461 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_16_), 
        .B0(n230), .B1(Input2[16]), .Y(n3228) );
  CLKINVX1 U3462 ( .A(n1013), .Y(n1012) );
  OAI2B2X1 U3463 ( .A1N(Input2[16]), .A0(n3153), .B0(n3229), .B1(n3152), .Y(
        n1013) );
  CLKINVX1 U3464 ( .A(Output2[16]), .Y(n3229) );
  XOR2X1 U3465 ( .A(n3230), .B(n1256), .Y(Output2[16]) );
  AOI221XL U3466 ( .A0(n3160), .A1(n296), .B0(n3182), .B1(n2293), .C0(n3231), 
        .Y(n1256) );
  AO22X1 U3467 ( .A0(n266), .A1(n3232), .B0(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]), .B1(n292), .Y(n3231) );
  CLKINVX1 U3468 ( .A(n2011), .Y(n3182) );
  MXI2X1 U3469 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .B(n3233), .S0(
        n310), .Y(n2011) );
  XOR2X1 U3470 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[25]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[121]), .Y(n3233) );
  XOR2X1 U3471 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_4_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]), .Y(n3160) );
  CLKNAND2X2 U3472 ( .A(Input2[16]), .B(n2288), .Y(n3230) );
  OAI221X1 U3473 ( .A0(n3234), .A1(n2300), .B0(n3235), .B1(n2302), .C0(n3236), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_15_N3) );
  AOI22XL U3474 ( .A0(n186), .A1(n1016), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1258), .Y(n3236) );
  OAI2B2X1 U3475 ( .A1N(Output2[15]), .A0(n2379), .B0(n3235), .B1(n2381), .Y(
        n1016) );
  XOR2X1 U3476 ( .A(n1258), .B(n3237), .Y(Output2[15]) );
  NOR2X1 U3477 ( .A(n248), .B(n3235), .Y(n3237) );
  OAI221X1 U3478 ( .A0(n2020), .A1(n277), .B0(n2267), .B1(n3238), .C0(n3239), 
        .Y(n1258) );
  AOI222XL U3479 ( .A0(n260), .A1(n3240), .B0(n2258), .B1(n3241), .C0(n2312), 
        .C1(n2499), .Y(n3239) );
  XOR2X1 U3480 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_2_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[23]), .Y(n2499) );
  XOR2X1 U3481 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[112]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]), .Y(n3241) );
  CLKINVX1 U3482 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .Y(n3238) );
  CLKINVX1 U3483 ( .A(Input2[15]), .Y(n3235) );
  CLKINVX1 U3484 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_15_), .Y(n3234) );
  OAI221X1 U3485 ( .A0(n1019), .A1(n175), .B0(n1259), .B1(n147), .C0(n3242), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_14_N3) );
  AOI22XL U3486 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_14_), 
        .B0(n229), .B1(Input2[14]), .Y(n3242) );
  CLKINVX1 U3487 ( .A(n1020), .Y(n1019) );
  OAI2B2X1 U3488 ( .A1N(Output2[14]), .A0(n2379), .B0(n3243), .B1(n2381), .Y(
        n1020) );
  CLKINVX1 U3489 ( .A(Input2[14]), .Y(n3243) );
  XOR2X1 U3490 ( .A(n3244), .B(n1259), .Y(Output2[14]) );
  CLKINVX1 U3491 ( .A(n3245), .Y(n1259) );
  OAI221X1 U3492 ( .A0(n3246), .A1(n2274), .B0(n3247), .B1(n2273), .C0(n3248), 
        .Y(n3245) );
  AOI22XL U3493 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[10]), .A1(n297), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .B1(n292), .Y(n3248) );
  XOR2X1 U3494 ( .A(n3249), .B(n3250), .Y(n3246) );
  MXI2X1 U3495 ( .A(n2724), .B(n3251), .S0(n310), .Y(n3250) );
  XOR2X1 U3496 ( .A(n3252), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[20]), .Y(
        n3251) );
  CLKINVX1 U3497 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[12]), .Y(n2724) );
  OR2X1 U3498 ( .A(n2015), .B(n2133), .Y(n3249) );
  MXI2X1 U3499 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[15]), .B(n3253), .S0(
        n310), .Y(n2133) );
  XOR2X1 U3500 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[23]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[119]), .Y(n3253) );
  CLKNAND2X2 U3501 ( .A(Input2[14]), .B(n2288), .Y(n3244) );
  OAI221X1 U3502 ( .A0(n1023), .A1(n175), .B0(n3254), .B1(n147), .C0(n3255), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_13_N3) );
  AOI22XL U3503 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_13_), 
        .B0(n229), .B1(Input2[13]), .Y(n3255) );
  CLKINVX1 U3504 ( .A(n1261), .Y(n3254) );
  CLKINVX1 U3505 ( .A(n1024), .Y(n1023) );
  OAI2B2X1 U3506 ( .A1N(Output2[13]), .A0(n2379), .B0(n3256), .B1(n2381), .Y(
        n1024) );
  XOR2X1 U3507 ( .A(n1261), .B(n3257), .Y(Output2[13]) );
  NOR2X1 U3508 ( .A(n248), .B(n3256), .Y(n3257) );
  CLKINVX1 U3509 ( .A(Input2[13]), .Y(n3256) );
  OAI222X1 U3510 ( .A0(n2730), .A1(n2135), .B0(n3258), .B1(n2274), .C0(n3259), 
        .C1(n2273), .Y(n1261) );
  XOR2X1 U3511 ( .A(n3260), .B(n3261), .Y(n3258) );
  MXI2X1 U3512 ( .A(n3262), .B(n3263), .S0(n310), .Y(n3261) );
  XOR2X1 U3513 ( .A(n3264), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[16]), .Y(
        n3263) );
  CLKINVX1 U3514 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[8]), .Y(n3262) );
  CLKNAND2X2 U3515 ( .A(n3265), .B(n2500), .Y(n3260) );
  CLKINVX1 U3516 ( .A(n2018), .Y(n2500) );
  MXI2X1 U3517 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .B(n3266), .S0(
        n310), .Y(n2018) );
  XOR2X1 U3518 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[113]), .Y(n3266) );
  OAI221X1 U3519 ( .A0(n3267), .A1(n2300), .B0(n3268), .B1(n2302), .C0(n3269), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_127_N3) );
  AOI22XL U3520 ( .A0(n186), .A1(n589), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1072), .Y(n3269) );
  CLKINVX1 U3521 ( .A(n586), .Y(n589) );
  MXI2X1 U3522 ( .A(Input2[127]), .B(Output2[127]), .S0(dec), .Y(n586) );
  XOR2X1 U3523 ( .A(n1072), .B(n3270), .Y(Output2[127]) );
  NOR2X1 U3524 ( .A(n248), .B(n3268), .Y(n3270) );
  OAI221X1 U3525 ( .A0(n2032), .A1(n278), .B0(n2267), .B1(n3271), .C0(n3272), 
        .Y(n1072) );
  AOI222XL U3526 ( .A0(n2312), .A1(n3273), .B0(n2258), .B1(n3274), .C0(n265), 
        .C1(n3275), .Y(n3272) );
  XNOR2X1 U3527 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[31]), .B(n3071), .Y(
        n3275) );
  XNOR2X1 U3528 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[63]), .B(n2307), .Y(
        n3071) );
  XOR2X1 U3529 ( .A(n3276), .B(n3277), .Y(n2307) );
  XOR2X1 U3530 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[88]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_53_), .Y(n3274) );
  CLKINVX1 U3531 ( .A(Input2[127]), .Y(n3268) );
  CLKINVX1 U3532 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_127_), .Y(n3267) );
  OAI221X1 U3533 ( .A0(n592), .A1(n175), .B0(n1073), .B1(n147), .C0(n3278), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_126_N3) );
  AOI22XL U3534 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_126_), 
        .B0(n229), .B1(Input2[126]), .Y(n3278) );
  MXI2X1 U3535 ( .A(Input2[126]), .B(Output2[126]), .S0(dec), .Y(n592) );
  XOR2X1 U3536 ( .A(n3279), .B(n1073), .Y(Output2[126]) );
  CLKINVX1 U3537 ( .A(n3280), .Y(n1073) );
  OAI221X1 U3538 ( .A0(n3281), .A1(n2273), .B0(n3282), .B1(n2274), .C0(n3283), 
        .Y(n3280) );
  AOI22XL U3539 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[122]), .A1(n298), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[121]), .B1(n292), .Y(n3283) );
  XOR2X1 U3540 ( .A(n3284), .B(n3285), .Y(n3282) );
  MXI2X1 U3541 ( .A(n3171), .B(n3286), .S0(n311), .Y(n3285) );
  XOR2X1 U3542 ( .A(n3287), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[92]), .Y(
        n3286) );
  OR2X1 U3543 ( .A(n2145), .B(n2026), .Y(n3284) );
  XOR2X1 U3544 ( .A(n3081), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[20]), .Y(
        n3281) );
  XOR2X1 U3545 ( .A(n2913), .B(n2320), .Y(n3081) );
  XOR2X1 U3546 ( .A(n3288), .B(n3171), .Y(n2320) );
  CLKINVX1 U3547 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[124]), .Y(n3171) );
  CLKINVX1 U3548 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[44]), .Y(n2913) );
  CLKNAND2X2 U3549 ( .A(Input2[126]), .B(n2288), .Y(n3279) );
  OAI221X1 U3550 ( .A0(n595), .A1(n175), .B0(n1074), .B1(n147), .C0(n3289), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_125_N3) );
  AOI22XL U3551 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_125_), 
        .B0(n229), .B1(Input2[125]), .Y(n3289) );
  MXI2X1 U3552 ( .A(Input2[125]), .B(Output2[125]), .S0(dec), .Y(n595) );
  XOR2X1 U3553 ( .A(n3290), .B(n1074), .Y(Output2[125]) );
  CLKINVX1 U3554 ( .A(n3291), .Y(n1074) );
  OAI222X1 U3555 ( .A0(n3292), .A1(n2274), .B0(n3293), .B1(n2273), .C0(n2730), 
        .C1(n2147), .Y(n3291) );
  XOR2X1 U3556 ( .A(n3102), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[16]), .Y(
        n3293) );
  XOR2X1 U3557 ( .A(n2924), .B(n2334), .Y(n3102) );
  XNOR2X1 U3558 ( .A(n3294), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[120]), .Y(
        n2334) );
  CLKINVX1 U3559 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[40]), .Y(n2924) );
  XOR2X1 U3560 ( .A(n3295), .B(n3296), .Y(n3292) );
  MXI2X1 U3561 ( .A(n3181), .B(n3297), .S0(n311), .Y(n3296) );
  XOR2X1 U3562 ( .A(n3298), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[88]), .Y(
        n3297) );
  CLKINVX1 U3563 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[120]), .Y(n3181) );
  OR2X1 U3564 ( .A(n2030), .B(n2149), .Y(n3295) );
  CLKNAND2X2 U3565 ( .A(Input2[125]), .B(n2288), .Y(n3290) );
  OAI221X1 U3566 ( .A0(n598), .A1(n175), .B0(n3299), .B1(n147), .C0(n3300), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_124_N3) );
  AOI22XL U3567 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_124_), 
        .B0(n229), .B1(Input2[124]), .Y(n3300) );
  CLKINVX1 U3568 ( .A(n1076), .Y(n3299) );
  MXI2X1 U3569 ( .A(Input2[124]), .B(Output2[124]), .S0(dec), .Y(n598) );
  XOR2X1 U3570 ( .A(n1076), .B(n3301), .Y(Output2[124]) );
  NOR2BX1 U3571 ( .AN(Input2[124]), .B(n254), .Y(n3301) );
  OAI221X1 U3572 ( .A0(n2149), .A1(n2274), .B0(n276), .B1(n2028), .C0(n3302), 
        .Y(n1076) );
  AOI22XL U3573 ( .A0(n263), .A1(n3303), .B0(n295), .B1(n3304), .Y(n3302) );
  XNOR2X1 U3574 ( .A(n3113), .B(n2131), .Y(n3303) );
  XNOR2X1 U3575 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_5_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[19]), .Y(n2131) );
  XNOR2X1 U3576 ( .A(n2349), .B(n2232), .Y(n3113) );
  XNOR2X1 U3577 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_11_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[43]), .Y(n2232) );
  XOR2X1 U3578 ( .A(n3287), .B(n2151), .Y(n2349) );
  MXI2X1 U3579 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[123]), .B(n3305), .S0(
        n311), .Y(n2149) );
  XOR2X1 U3580 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[91]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_51_), .Y(n3305) );
  OAI221X1 U3581 ( .A0(n601), .A1(n175), .B0(n3306), .B1(n147), .C0(n3307), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_123_N3) );
  AOI22XL U3582 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_123_), 
        .B0(n229), .B1(Input2[123]), .Y(n3307) );
  CLKINVX1 U3583 ( .A(n1078), .Y(n3306) );
  MXI2X1 U3584 ( .A(Input2[123]), .B(Output2[123]), .S0(dec), .Y(n601) );
  XOR2X1 U3585 ( .A(n1078), .B(n3308), .Y(Output2[123]) );
  NOR2BX1 U3586 ( .AN(Input2[123]), .B(n255), .Y(n3308) );
  OAI211XL U3587 ( .A0(n2255), .A1(n3309), .B0(n3310), .C0(n3311), .Y(n1078)
         );
  AOI22XL U3588 ( .A0(n2258), .A1(n3312), .B0(n261), .B1(n3313), .Y(n3311) );
  XOR2X1 U3589 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[17]), .B(n3119), .Y(
        n3313) );
  XNOR2X1 U3590 ( .A(n2897), .B(n2357), .Y(n3119) );
  XOR2X1 U3591 ( .A(n3314), .B(n3271), .Y(n2357) );
  CLKINVX1 U3592 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[121]), .Y(n3271) );
  CLKINVX1 U3593 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[41]), .Y(n2897) );
  XOR2X1 U3594 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[90]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_50_), .Y(n3312) );
  MXI2X1 U3595 ( .A(n3315), .B(n3316), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[124]), .Y(n3310) );
  OAI21X1 U3596 ( .A0(n3317), .A1(n281), .B0(n2267), .Y(n3316) );
  NOR2X1 U3597 ( .A(n2028), .B(n2147), .Y(n3317) );
  NOR3X1 U3598 ( .A(n2147), .B(n276), .C(n2028), .Y(n3315) );
  CLKINVX1 U3599 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[127]), .Y(n2147) );
  OAI221X1 U3600 ( .A0(n604), .A1(n175), .B0(n3318), .B1(n147), .C0(n3319), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_122_N3) );
  AOI22XL U3601 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_122_), 
        .B0(n229), .B1(Input2[122]), .Y(n3319) );
  CLKINVX1 U3602 ( .A(n1080), .Y(n3318) );
  MXI2X1 U3603 ( .A(Input2[122]), .B(Output2[122]), .S0(dec), .Y(n604) );
  XOR2X1 U3604 ( .A(n1080), .B(n3320), .Y(Output2[122]) );
  NOR2BX1 U3605 ( .AN(Input2[122]), .B(n254), .Y(n3320) );
  OAI221X1 U3606 ( .A0(n3321), .A1(n2273), .B0(n2026), .B1(n2274), .C0(n3322), 
        .Y(n1080) );
  MXI2X1 U3607 ( .A(n3323), .B(n3324), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[120]), .Y(n3322) );
  OAI21X1 U3608 ( .A0(n3325), .A1(n281), .B0(n2267), .Y(n3324) );
  NOR2X1 U3609 ( .A(n2151), .B(n2032), .Y(n3325) );
  NOR3X1 U3610 ( .A(n282), .B(n2151), .C(n2032), .Y(n3323) );
  MXI2X1 U3611 ( .A(n3304), .B(n3326), .S0(n311), .Y(n2026) );
  XOR2X1 U3612 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[92]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_54_), .Y(n3326) );
  XNOR2X1 U3613 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_31_), .B(n2028), .Y(
        n3304) );
  CLKINVX1 U3614 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[124]), .Y(n2028) );
  XOR2X1 U3615 ( .A(n3130), .B(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]), .Y(
        n3321) );
  XOR2X1 U3616 ( .A(n2106), .B(n2370), .Y(n3130) );
  XNOR2X1 U3617 ( .A(n3327), .B(Inst_forkAE_CipherInst_RF_S_MID_C2[124]), .Y(
        n2370) );
  CLKINVX1 U3618 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[58]), .Y(n2106) );
  OAI221X1 U3619 ( .A0(n607), .A1(n175), .B0(n1081), .B1(n147), .C0(n3328), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_121_N3) );
  AOI22XL U3620 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_121_), 
        .B0(n229), .B1(Input2[121]), .Y(n3328) );
  MXI2X1 U3621 ( .A(Input2[121]), .B(Output2[121]), .S0(dec), .Y(n607) );
  XOR2X1 U3622 ( .A(n3329), .B(n1081), .Y(Output2[121]) );
  CLKINVX1 U3623 ( .A(n3330), .Y(n1081) );
  OAI221X1 U3624 ( .A0(n3331), .A1(n2273), .B0(n2145), .B1(n2274), .C0(n3332), 
        .Y(n3330) );
  AOI2BB2X1 U3625 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[123]), .B1(n294), 
        .A0N(n285), .A1N(n2151), .Y(n3332) );
  XNOR2X1 U3626 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_31_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[123]), .Y(n2151) );
  MXI2X1 U3627 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[127]), .B(n3333), .S0(
        n311), .Y(n2145) );
  XOR2X1 U3628 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[95]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_55_), .Y(n3333) );
  XOR2X1 U3629 ( .A(n3140), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[23]), .Y(
        n3331) );
  XOR2X1 U3630 ( .A(n2229), .B(n2392), .Y(n3140) );
  XOR2X1 U3631 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_49_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[127]), .Y(n2392) );
  CLKINVX1 U3632 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[47]), .Y(n2229) );
  CLKNAND2X2 U3633 ( .A(Input2[121]), .B(n2288), .Y(n3329) );
  OAI221X1 U3634 ( .A0(n610), .A1(n175), .B0(n3334), .B1(n147), .C0(n3335), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_120_N3) );
  AOI22XL U3635 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_120_), 
        .B0(n229), .B1(Input2[120]), .Y(n3335) );
  CLKINVX1 U3636 ( .A(n1083), .Y(n3334) );
  MXI2X1 U3637 ( .A(Input2[120]), .B(Output2[120]), .S0(dec), .Y(n610) );
  XOR2X1 U3638 ( .A(n1083), .B(n3336), .Y(Output2[120]) );
  NOR2BX1 U3639 ( .AN(Input2[120]), .B(n254), .Y(n3336) );
  OAI221X1 U3640 ( .A0(n2030), .A1(n2274), .B0(n275), .B1(n3277), .C0(n3337), 
        .Y(n1083) );
  AOI22XL U3641 ( .A0(n264), .A1(n3338), .B0(n295), .B1(n3273), .Y(n3337) );
  XNOR2X1 U3642 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_30_), .B(n3277), .Y(
        n3273) );
  XOR2X1 U3643 ( .A(n3147), .B(n3158), .Y(n3338) );
  CLKINVX1 U3644 ( .A(n2013), .Y(n3158) );
  XNOR2X1 U3645 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_4_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[18]), .Y(n2013) );
  XNOR2X1 U3646 ( .A(n2400), .B(n2109), .Y(n3147) );
  XNOR2X1 U3647 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_10_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[42]), .Y(n2109) );
  XOR2X1 U3648 ( .A(n3298), .B(n2032), .Y(n2400) );
  XOR2X1 U3649 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_30_), .B(n3309), .Y(
        n2032) );
  CLKINVX1 U3650 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[122]), .Y(n3309) );
  CLKINVX1 U3651 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[120]), .Y(n3277) );
  MXI2X1 U3652 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[121]), .B(n3339), .S0(
        n311), .Y(n2030) );
  XOR2X1 U3653 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[89]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_49_), .Y(n3339) );
  OAI221X1 U3654 ( .A0(n1027), .A1(n175), .B0(n1263), .B1(n147), .C0(n3340), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_12_N3) );
  AOI22XL U3655 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_12_), 
        .B0(n229), .B1(Input2[12]), .Y(n3340) );
  CLKINVX1 U3656 ( .A(n1028), .Y(n1027) );
  OAI2B2X1 U3657 ( .A1N(Input2[12]), .A0(n2381), .B0(n3341), .B1(n2379), .Y(
        n1028) );
  CLKINVX1 U3658 ( .A(Output2[12]), .Y(n3341) );
  XOR2X1 U3659 ( .A(n3342), .B(n1263), .Y(Output2[12]) );
  AOI221XL U3660 ( .A0(n3343), .A1(n296), .B0(n3265), .B1(n2293), .C0(n3344), 
        .Y(n1263) );
  OAI2BB2X1 U3661 ( .B0(n2017), .B1(n284), .A0N(n3345), .A1N(n268), .Y(n3344)
         );
  CLKINVX1 U3662 ( .A(n2137), .Y(n3265) );
  MXI2X1 U3663 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[11]), .B(n3346), .S0(
        n311), .Y(n2137) );
  XOR2X1 U3664 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[19]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[115]), .Y(n3346) );
  CLKNAND2X2 U3665 ( .A(Input2[12]), .B(n2288), .Y(n3342) );
  OAI221X1 U3666 ( .A0(n3347), .A1(n2300), .B0(n3348), .B1(n2302), .C0(n3349), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_119_N3) );
  AOI22XL U3667 ( .A0(n186), .A1(n613), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1085), .Y(n3349) );
  OAI2B2X1 U3668 ( .A1N(Output2[119]), .A0(n3350), .B0(n3348), .B1(n3351), .Y(
        n613) );
  XOR2X1 U3669 ( .A(n1085), .B(n3352), .Y(Output2[119]) );
  NOR2X1 U3670 ( .A(n248), .B(n3348), .Y(n3352) );
  OAI221X1 U3671 ( .A0(n2040), .A1(n278), .B0(n2267), .B1(n3353), .C0(n3354), 
        .Y(n1085) );
  AOI222XL U3672 ( .A0(n2312), .A1(n3355), .B0(n2258), .B1(n3356), .C0(n264), 
        .C1(n3357), .Y(n3354) );
  XOR2X1 U3673 ( .A(n2502), .B(n3155), .Y(n3357) );
  XOR2X1 U3674 ( .A(n3060), .B(n2410), .Y(n3155) );
  XOR2X1 U3675 ( .A(n3358), .B(n3359), .Y(n2410) );
  CLKINVX1 U3676 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[55]), .Y(n3060) );
  CLKINVX1 U3677 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[23]), .Y(n2502) );
  XOR2X1 U3678 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[80]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_5_), .Y(n3356) );
  CLKINVX1 U3679 ( .A(Input2[119]), .Y(n3348) );
  CLKINVX1 U3680 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_119_), .Y(n3347) );
  OAI221X1 U3681 ( .A0(n616), .A1(n175), .B0(n1086), .B1(n147), .C0(n3360), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_118_N3) );
  AOI22XL U3682 ( .A0(n201), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_118_), 
        .B0(n229), .B1(Input2[118]), .Y(n3360) );
  CLKINVX1 U3683 ( .A(n617), .Y(n616) );
  OAI2B2X1 U3684 ( .A1N(Output2[118]), .A0(n3350), .B0(n3361), .B1(n3351), .Y(
        n617) );
  CLKINVX1 U3685 ( .A(Input2[118]), .Y(n3361) );
  XOR2X1 U3686 ( .A(n3362), .B(n1086), .Y(Output2[118]) );
  CLKINVX1 U3687 ( .A(n3363), .Y(n1086) );
  OAI221X1 U3688 ( .A0(n3364), .A1(n2273), .B0(n3365), .B1(n2274), .C0(n3366), 
        .Y(n3363) );
  AOI22XL U3689 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[114]), .A1(n298), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[113]), .B1(n292), .Y(n3366) );
  XOR2X1 U3690 ( .A(n3367), .B(n3368), .Y(n3365) );
  MXI2X1 U3691 ( .A(n3252), .B(n3369), .S0(n311), .Y(n3368) );
  XOR2X1 U3692 ( .A(n3370), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[84]), .Y(
        n3369) );
  OR2X1 U3693 ( .A(n2153), .B(n2034), .Y(n3367) );
  XOR2X1 U3694 ( .A(n3166), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[12]), .Y(
        n3364) );
  XOR2X1 U3695 ( .A(n3003), .B(n2422), .Y(n3166) );
  XOR2X1 U3696 ( .A(n3371), .B(n3252), .Y(n2422) );
  CLKINVX1 U3697 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[116]), .Y(n3252) );
  CLKINVX1 U3698 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[36]), .Y(n3003) );
  CLKNAND2X2 U3699 ( .A(Input2[118]), .B(n2288), .Y(n3362) );
  OAI221X1 U3700 ( .A0(n620), .A1(n174), .B0(n1087), .B1(n146), .C0(n3372), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_117_N3) );
  AOI22XL U3701 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_117_), 
        .B0(n229), .B1(Input2[117]), .Y(n3372) );
  CLKINVX1 U3702 ( .A(n621), .Y(n620) );
  OAI2B2X1 U3703 ( .A1N(Output2[117]), .A0(n3350), .B0(n3373), .B1(n3351), .Y(
        n621) );
  CLKINVX1 U3704 ( .A(Input2[117]), .Y(n3373) );
  XOR2X1 U3705 ( .A(n3374), .B(n1087), .Y(Output2[117]) );
  CLKINVX1 U3706 ( .A(n3375), .Y(n1087) );
  OAI222X1 U3707 ( .A0(n3376), .A1(n2274), .B0(n3377), .B1(n2273), .C0(n2730), 
        .C1(n2155), .Y(n3375) );
  XOR2X1 U3708 ( .A(n3177), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[8]), .Y(
        n3377) );
  XOR2X1 U3709 ( .A(n3014), .B(n2435), .Y(n3177) );
  XNOR2X1 U3710 ( .A(n3378), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[112]), .Y(
        n2435) );
  CLKINVX1 U3711 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[32]), .Y(n3014) );
  XOR2X1 U3712 ( .A(n3379), .B(n3380), .Y(n3376) );
  MXI2X1 U3713 ( .A(n3264), .B(n3381), .S0(n311), .Y(n3380) );
  XOR2X1 U3714 ( .A(n3382), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[80]), .Y(
        n3381) );
  CLKINVX1 U3715 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[112]), .Y(n3264) );
  OR2X1 U3716 ( .A(n2038), .B(n2157), .Y(n3379) );
  CLKNAND2X2 U3717 ( .A(Input2[117]), .B(n2288), .Y(n3374) );
  OAI221X1 U3718 ( .A0(n624), .A1(n174), .B0(n3383), .B1(n146), .C0(n3384), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_116_N3) );
  AOI22XL U3719 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_116_), 
        .B0(n229), .B1(Input2[116]), .Y(n3384) );
  CLKINVX1 U3720 ( .A(n1089), .Y(n3383) );
  CLKINVX1 U3721 ( .A(n625), .Y(n624) );
  OAI2B2X1 U3722 ( .A1N(Output2[116]), .A0(n3350), .B0(n3385), .B1(n3351), .Y(
        n625) );
  XOR2X1 U3723 ( .A(n1089), .B(n3386), .Y(Output2[116]) );
  NOR2X1 U3724 ( .A(n248), .B(n3385), .Y(n3386) );
  CLKINVX1 U3725 ( .A(Input2[116]), .Y(n3385) );
  OAI221X1 U3726 ( .A0(n2157), .A1(n2274), .B0(n274), .B1(n2036), .C0(n3387), 
        .Y(n1089) );
  AOI22XL U3727 ( .A0(n262), .A1(n3388), .B0(n295), .B1(n3389), .Y(n3387) );
  XOR2X1 U3728 ( .A(n2386), .B(n3189), .Y(n3388) );
  XNOR2X1 U3729 ( .A(n2450), .B(n2239), .Y(n3189) );
  XNOR2X1 U3730 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_9_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[35]), .Y(n2239) );
  XOR2X1 U3731 ( .A(n3370), .B(n2159), .Y(n2450) );
  MXI2X1 U3732 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[115]), .B(n3390), .S0(
        n311), .Y(n2157) );
  XOR2X1 U3733 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[83]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_3_), .Y(n3390) );
  OAI221X1 U3734 ( .A0(n628), .A1(n174), .B0(n3391), .B1(n146), .C0(n3392), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_115_N3) );
  AOI22XL U3735 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_115_), 
        .B0(n228), .B1(Input2[115]), .Y(n3392) );
  CLKINVX1 U3736 ( .A(n1091), .Y(n3391) );
  CLKINVX1 U3737 ( .A(n629), .Y(n628) );
  OAI2B2X1 U3738 ( .A1N(Output2[115]), .A0(n3350), .B0(n3393), .B1(n3351), .Y(
        n629) );
  XOR2X1 U3739 ( .A(n1091), .B(n3394), .Y(Output2[115]) );
  NOR2X1 U3740 ( .A(n248), .B(n3393), .Y(n3394) );
  CLKINVX1 U3741 ( .A(Input2[115]), .Y(n3393) );
  OAI211XL U3742 ( .A0(n2255), .A1(n3395), .B0(n3396), .C0(n3397), .Y(n1091)
         );
  AOI22XL U3743 ( .A0(n2258), .A1(n3398), .B0(n261), .B1(n3399), .Y(n3397) );
  XOR2X1 U3744 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .B(n3204), .Y(
        n3399) );
  XNOR2X1 U3745 ( .A(n2987), .B(n2458), .Y(n3204) );
  XOR2X1 U3746 ( .A(n3400), .B(n3353), .Y(n2458) );
  CLKINVX1 U3747 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[113]), .Y(n3353) );
  CLKINVX1 U3748 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[33]), .Y(n2987) );
  XOR2X1 U3749 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[82]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_2_), .Y(n3398) );
  MXI2X1 U3750 ( .A(n3401), .B(n3402), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[116]), .Y(n3396) );
  OAI21X1 U3751 ( .A0(n3403), .A1(n281), .B0(n2267), .Y(n3402) );
  NOR2X1 U3752 ( .A(n2155), .B(n2036), .Y(n3403) );
  NOR3X1 U3753 ( .A(n2036), .B(n2155), .C(n278), .Y(n3401) );
  CLKINVX1 U3754 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[119]), .Y(n2155) );
  OAI221X1 U3755 ( .A0(n632), .A1(n174), .B0(n3404), .B1(n146), .C0(n3405), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_114_N3) );
  AOI22XL U3756 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_114_), 
        .B0(n228), .B1(Input2[114]), .Y(n3405) );
  CLKINVX1 U3757 ( .A(n1093), .Y(n3404) );
  CLKINVX1 U3758 ( .A(n633), .Y(n632) );
  OAI2B2X1 U3759 ( .A1N(Output2[114]), .A0(n3350), .B0(n3406), .B1(n3351), .Y(
        n633) );
  XOR2X1 U3760 ( .A(n1093), .B(n3407), .Y(Output2[114]) );
  NOR2X1 U3761 ( .A(n248), .B(n3406), .Y(n3407) );
  CLKINVX1 U3762 ( .A(Input2[114]), .Y(n3406) );
  OAI221X1 U3763 ( .A0(n3408), .A1(n2273), .B0(n2034), .B1(n2274), .C0(n3409), 
        .Y(n1093) );
  MXI2X1 U3764 ( .A(n3410), .B(n3411), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[112]), .Y(n3409) );
  OAI21X1 U3765 ( .A0(n3412), .A1(n281), .B0(n2267), .Y(n3411) );
  NOR2X1 U3766 ( .A(n2159), .B(n2040), .Y(n3412) );
  NOR3X1 U3767 ( .A(n274), .B(n2159), .C(n2040), .Y(n3410) );
  MXI2X1 U3768 ( .A(n3389), .B(n3413), .S0(n311), .Y(n2034) );
  XOR2X1 U3769 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[84]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_6_), .Y(n3413) );
  XNOR2X1 U3770 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_29_), .B(n2036), .Y(
        n3389) );
  CLKINVX1 U3771 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[116]), .Y(n2036) );
  XOR2X1 U3772 ( .A(n3215), .B(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]), .Y(
        n3408) );
  XOR2X1 U3773 ( .A(n2113), .B(n2471), .Y(n3215) );
  XNOR2X1 U3774 ( .A(n3414), .B(Inst_forkAE_CipherInst_RF_S_MID_C2[116]), .Y(
        n2471) );
  CLKINVX1 U3775 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[50]), .Y(n2113) );
  OAI221X1 U3776 ( .A0(n636), .A1(n174), .B0(n1094), .B1(n146), .C0(n3415), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_113_N3) );
  AOI22XL U3777 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_113_), 
        .B0(n228), .B1(Input2[113]), .Y(n3415) );
  CLKINVX1 U3778 ( .A(n637), .Y(n636) );
  OAI2B2X1 U3779 ( .A1N(Output2[113]), .A0(n3350), .B0(n3416), .B1(n3351), .Y(
        n637) );
  CLKINVX1 U3780 ( .A(Input2[113]), .Y(n3416) );
  XOR2X1 U3781 ( .A(n3417), .B(n1094), .Y(Output2[113]) );
  CLKINVX1 U3782 ( .A(n3418), .Y(n1094) );
  OAI221X1 U3783 ( .A0(n3419), .A1(n2273), .B0(n2153), .B1(n2274), .C0(n3420), 
        .Y(n3418) );
  AOI2BB2X1 U3784 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[115]), .B1(n294), 
        .A0N(n285), .A1N(n2159), .Y(n3420) );
  XNOR2X1 U3785 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_29_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[115]), .Y(n2159) );
  MXI2X1 U3786 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[119]), .B(n3421), .S0(
        n311), .Y(n2153) );
  XOR2X1 U3787 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[87]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_7_), .Y(n3421) );
  XOR2X1 U3788 ( .A(n3226), .B(n2135), .Y(n3419) );
  XNOR2X1 U3789 ( .A(n2236), .B(n2484), .Y(n3226) );
  XOR2X1 U3790 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_1_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[119]), .Y(n2484) );
  CLKINVX1 U3791 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[39]), .Y(n2236) );
  CLKNAND2X2 U3792 ( .A(Input2[113]), .B(n2288), .Y(n3417) );
  OAI221X1 U3793 ( .A0(n640), .A1(n174), .B0(n3422), .B1(n146), .C0(n3423), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_112_N3) );
  AOI22XL U3794 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_112_), 
        .B0(n228), .B1(Input2[112]), .Y(n3423) );
  CLKINVX1 U3795 ( .A(n1096), .Y(n3422) );
  CLKINVX1 U3796 ( .A(n641), .Y(n640) );
  OAI2B2X1 U3797 ( .A1N(Output2[112]), .A0(n3350), .B0(n3424), .B1(n3351), .Y(
        n641) );
  XOR2X1 U3798 ( .A(n1096), .B(n3425), .Y(Output2[112]) );
  NOR2X1 U3799 ( .A(n249), .B(n3424), .Y(n3425) );
  CLKINVX1 U3800 ( .A(Input2[112]), .Y(n3424) );
  OAI221X1 U3801 ( .A0(n2038), .A1(n2274), .B0(n281), .B1(n3359), .C0(n3426), 
        .Y(n1096) );
  AOI22XL U3802 ( .A0(n263), .A1(n3427), .B0(n295), .B1(n3355), .Y(n3426) );
  XNOR2X1 U3803 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_28_), .B(n3359), .Y(
        n3355) );
  XNOR2X1 U3804 ( .A(n3232), .B(n2020), .Y(n3427) );
  XNOR2X1 U3805 ( .A(n2492), .B(n2116), .Y(n3232) );
  XNOR2X1 U3806 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_8_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[34]), .Y(n2116) );
  XOR2X1 U3807 ( .A(n3382), .B(n2040), .Y(n2492) );
  XOR2X1 U3808 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_28_), .B(n3395), .Y(
        n2040) );
  CLKINVX1 U3809 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[114]), .Y(n3395) );
  CLKINVX1 U3810 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[112]), .Y(n3359) );
  MXI2X1 U3811 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[113]), .B(n3428), .S0(
        n316), .Y(n2038) );
  XOR2X1 U3812 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[81]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_1_), .Y(n3428) );
  OAI221X1 U3813 ( .A0(n3429), .A1(n2300), .B0(n3430), .B1(n2302), .C0(n3431), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_111_N3) );
  AOI22XL U3814 ( .A0(n186), .A1(n644), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1098), .Y(n3431) );
  OAI2B2X1 U3815 ( .A1N(Output2[111]), .A0(n3432), .B0(n3430), .B1(n3433), .Y(
        n644) );
  XOR2X1 U3816 ( .A(n1098), .B(n3434), .Y(Output2[111]) );
  NOR2X1 U3817 ( .A(n249), .B(n3430), .Y(n3434) );
  OAI221X1 U3818 ( .A0(n2052), .A1(n277), .B0(n2267), .B1(n3435), .C0(n3436), 
        .Y(n1098) );
  AOI222XL U3819 ( .A0(n2312), .A1(n3437), .B0(n2258), .B1(n3438), .C0(n264), 
        .C1(n3439), .Y(n3436) );
  XOR2X1 U3820 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]), .B(n3240), .Y(
        n3439) );
  XOR2X1 U3821 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[47]), .B(n2518), .Y(
        n3240) );
  XNOR2X1 U3822 ( .A(n3440), .B(Inst_forkAE_CipherInst_RF_S_MID_C2[104]), .Y(
        n2518) );
  XOR2X1 U3823 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[72]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_61_), .Y(n3438) );
  CLKINVX1 U3824 ( .A(Input2[111]), .Y(n3430) );
  CLKINVX1 U3825 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_111_), .Y(n3429) );
  OAI221X1 U3826 ( .A0(n647), .A1(n174), .B0(n1099), .B1(n146), .C0(n3441), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_110_N3) );
  AOI22XL U3827 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_110_), 
        .B0(n228), .B1(Input2[110]), .Y(n3441) );
  CLKINVX1 U3828 ( .A(n648), .Y(n647) );
  OAI2B2X1 U3829 ( .A1N(Output2[110]), .A0(n3432), .B0(n3442), .B1(n3433), .Y(
        n648) );
  CLKINVX1 U3830 ( .A(Input2[110]), .Y(n3442) );
  XOR2X1 U3831 ( .A(n3443), .B(n1099), .Y(Output2[110]) );
  CLKINVX1 U3832 ( .A(n3444), .Y(n1099) );
  OAI221X1 U3833 ( .A0(n3445), .A1(n2273), .B0(n3446), .B1(n2274), .C0(n3447), 
        .Y(n3444) );
  AOI22XL U3834 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[106]), .A1(n298), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[105]), .B1(n291), .Y(n3447) );
  XOR2X1 U3835 ( .A(n3448), .B(n3449), .Y(n3446) );
  MXI2X1 U3836 ( .A(n2757), .B(n3450), .S0(n313), .Y(n3449) );
  XOR2X1 U3837 ( .A(n3451), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[76]), .Y(
        n3450) );
  OR2X1 U3838 ( .A(n2161), .B(n2042), .Y(n3448) );
  XOR2X1 U3839 ( .A(n3247), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[4]), .Y(
        n3445) );
  XOR2X1 U3840 ( .A(n2723), .B(n2523), .Y(n3247) );
  XOR2X1 U3841 ( .A(n3452), .B(n2757), .Y(n2523) );
  CLKINVX1 U3842 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[108]), .Y(n2757) );
  CLKINVX1 U3843 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[60]), .Y(n2723) );
  CLKNAND2X2 U3844 ( .A(Input2[110]), .B(n2288), .Y(n3443) );
  OAI221X1 U3845 ( .A0(n1031), .A1(n174), .B0(n3453), .B1(n146), .C0(n3454), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_11_N3) );
  AOI22XL U3846 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_11_), 
        .B0(n228), .B1(Input2[11]), .Y(n3454) );
  CLKINVX1 U3847 ( .A(n1265), .Y(n3453) );
  CLKINVX1 U3848 ( .A(n1032), .Y(n1031) );
  OAI2B2X1 U3849 ( .A1N(Output2[11]), .A0(n2379), .B0(n3455), .B1(n2381), .Y(
        n1032) );
  XOR2X1 U3850 ( .A(n1265), .B(n3456), .Y(Output2[11]) );
  NOR2X1 U3851 ( .A(n249), .B(n3455), .Y(n3456) );
  CLKINVX1 U3852 ( .A(Input2[11]), .Y(n3455) );
  OAI2B11X1 U3853 ( .A1N(n3457), .A0(n2273), .B0(n3458), .C0(n3459), .Y(n1265)
         );
  AOI22XL U3854 ( .A0(n2258), .A1(n3460), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[10]), .B1(n2312), .Y(n3459) );
  XOR2X1 U3855 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[18]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[114]), .Y(n3460) );
  MXI2X1 U3856 ( .A(n3461), .B(n3462), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[12]), .Y(n3458) );
  OAI21X1 U3857 ( .A0(n3463), .A1(n280), .B0(n2267), .Y(n3462) );
  NOR2X1 U3858 ( .A(n2135), .B(n2017), .Y(n3463) );
  NOR3X1 U3859 ( .A(n2017), .B(n2135), .C(n278), .Y(n3461) );
  CLKINVX1 U3860 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[15]), .Y(n2135) );
  CLKINVX1 U3861 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]), .Y(n2017) );
  OAI221X1 U3862 ( .A0(n651), .A1(n174), .B0(n1100), .B1(n146), .C0(n3464), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_109_N3) );
  AOI22XL U3863 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_109_), 
        .B0(n228), .B1(Input2[109]), .Y(n3464) );
  CLKINVX1 U3864 ( .A(n652), .Y(n651) );
  OAI2B2X1 U3865 ( .A1N(Output2[109]), .A0(n3432), .B0(n3465), .B1(n3433), .Y(
        n652) );
  CLKINVX1 U3866 ( .A(Input2[109]), .Y(n3465) );
  XOR2X1 U3867 ( .A(n3466), .B(n1100), .Y(Output2[109]) );
  CLKINVX1 U3868 ( .A(n3467), .Y(n1100) );
  OAI222X1 U3869 ( .A0(n3468), .A1(n2274), .B0(n3469), .B1(n2273), .C0(n2730), 
        .C1(n2163), .Y(n3467) );
  XOR2X1 U3870 ( .A(n3259), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[0]), .Y(
        n3469) );
  XOR2X1 U3871 ( .A(n2735), .B(n2536), .Y(n3259) );
  XNOR2X1 U3872 ( .A(n3470), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[104]), .Y(
        n2536) );
  CLKINVX1 U3873 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[56]), .Y(n2735) );
  XOR2X1 U3874 ( .A(n3471), .B(n3472), .Y(n3468) );
  MXI2X1 U3875 ( .A(n2871), .B(n3473), .S0(n312), .Y(n3472) );
  XOR2X1 U3876 ( .A(n3474), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[72]), .Y(
        n3473) );
  CLKINVX1 U3877 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[104]), .Y(n2871) );
  OR2X1 U3878 ( .A(n2050), .B(n2169), .Y(n3471) );
  CLKNAND2X2 U3879 ( .A(Input2[109]), .B(n2288), .Y(n3466) );
  OAI221X1 U3880 ( .A0(n655), .A1(n174), .B0(n3475), .B1(n146), .C0(n3476), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_108_N3) );
  AOI22XL U3881 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_108_), 
        .B0(n228), .B1(Input2[108]), .Y(n3476) );
  CLKINVX1 U3882 ( .A(n1102), .Y(n3475) );
  CLKINVX1 U3883 ( .A(n656), .Y(n655) );
  OAI2B2X1 U3884 ( .A1N(Output2[108]), .A0(n3432), .B0(n3477), .B1(n3433), .Y(
        n656) );
  XOR2X1 U3885 ( .A(n1102), .B(n3478), .Y(Output2[108]) );
  NOR2X1 U3886 ( .A(n249), .B(n3477), .Y(n3478) );
  CLKINVX1 U3887 ( .A(Input2[108]), .Y(n3477) );
  OAI221X1 U3888 ( .A0(n2169), .A1(n2274), .B0(n277), .B1(n2044), .C0(n3479), 
        .Y(n1102) );
  AOI22XL U3889 ( .A0(n263), .A1(n3480), .B0(n295), .B1(n3481), .Y(n3479) );
  XNOR2X1 U3890 ( .A(n2167), .B(n3345), .Y(n3480) );
  XNOR2X1 U3891 ( .A(n2551), .B(n2218), .Y(n3345) );
  XNOR2X1 U3892 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_15_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[59]), .Y(n2218) );
  XOR2X1 U3893 ( .A(n3451), .B(n2171), .Y(n2551) );
  MXI2X1 U3894 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[107]), .B(n3482), .S0(
        n310), .Y(n2169) );
  XOR2X1 U3895 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[75]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_59_), .Y(n3482) );
  OAI221X1 U3896 ( .A0(n659), .A1(n174), .B0(n3483), .B1(n146), .C0(n3484), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_107_N3) );
  AOI22XL U3897 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_107_), 
        .B0(n228), .B1(Input2[107]), .Y(n3484) );
  CLKINVX1 U3898 ( .A(n1104), .Y(n3483) );
  CLKINVX1 U3899 ( .A(n660), .Y(n659) );
  OAI2B2X1 U3900 ( .A1N(Output2[107]), .A0(n3432), .B0(n3485), .B1(n3433), .Y(
        n660) );
  XOR2X1 U3901 ( .A(n1104), .B(n3486), .Y(Output2[107]) );
  NOR2X1 U3902 ( .A(n249), .B(n3485), .Y(n3486) );
  CLKINVX1 U3903 ( .A(Input2[107]), .Y(n3485) );
  OAI211XL U3904 ( .A0(n2255), .A1(n3487), .B0(n3488), .C0(n3489), .Y(n1104)
         );
  AOI22XL U3905 ( .A0(n2258), .A1(n3490), .B0(n261), .B1(n3491), .Y(n3489) );
  XOR2X1 U3906 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .B(n3457), .Y(
        n3491) );
  XNOR2X1 U3907 ( .A(n2706), .B(n2559), .Y(n3457) );
  XOR2X1 U3908 ( .A(n3492), .B(n3435), .Y(n2559) );
  CLKINVX1 U3909 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[105]), .Y(n3435) );
  CLKINVX1 U3910 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[57]), .Y(n2706) );
  XOR2X1 U3911 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[74]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_58_), .Y(n3490) );
  MXI2X1 U3912 ( .A(n3493), .B(n3494), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[108]), .Y(n3488) );
  OAI21X1 U3913 ( .A0(n3495), .A1(n281), .B0(n2267), .Y(n3494) );
  NOR2X1 U3914 ( .A(n2163), .B(n2044), .Y(n3495) );
  NOR3X1 U3915 ( .A(n2044), .B(n2163), .C(n278), .Y(n3493) );
  CLKINVX1 U3916 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[111]), .Y(n2163) );
  OAI221X1 U3917 ( .A0(n663), .A1(n174), .B0(n3496), .B1(n146), .C0(n3497), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_106_N3) );
  AOI22XL U3918 ( .A0(n200), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_106_), 
        .B0(n228), .B1(Input2[106]), .Y(n3497) );
  CLKINVX1 U3919 ( .A(n1106), .Y(n3496) );
  CLKINVX1 U3920 ( .A(n664), .Y(n663) );
  OAI2B2X1 U3921 ( .A1N(Output2[106]), .A0(n3432), .B0(n3498), .B1(n3433), .Y(
        n664) );
  XOR2X1 U3922 ( .A(n1106), .B(n3499), .Y(Output2[106]) );
  NOR2X1 U3923 ( .A(n249), .B(n3498), .Y(n3499) );
  CLKINVX1 U3924 ( .A(Input2[106]), .Y(n3498) );
  OAI221X1 U3925 ( .A0(n3500), .A1(n2273), .B0(n2042), .B1(n2274), .C0(n3501), 
        .Y(n1106) );
  MXI2X1 U3926 ( .A(n3502), .B(n3503), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[104]), .Y(n3501) );
  OAI21X1 U3927 ( .A0(n3504), .A1(n281), .B0(n2267), .Y(n3503) );
  NOR2X1 U3928 ( .A(n2052), .B(n2171), .Y(n3504) );
  NOR3X1 U3929 ( .A(n274), .B(n2052), .C(n2171), .Y(n3502) );
  MXI2X1 U3930 ( .A(n3481), .B(n3505), .S0(n306), .Y(n2042) );
  XOR2X1 U3931 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[76]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_62_), .Y(n3505) );
  XNOR2X1 U3932 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_27_), .B(n2044), .Y(
        n3481) );
  CLKINVX1 U3933 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[108]), .Y(n2044) );
  XOR2X1 U3934 ( .A(n3506), .B(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[10]), .Y(
        n3500) );
  OAI221X1 U3935 ( .A0(n667), .A1(n173), .B0(n1107), .B1(n146), .C0(n3507), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_105_N3) );
  AOI22XL U3936 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_105_), 
        .B0(n228), .B1(Input2[105]), .Y(n3507) );
  CLKINVX1 U3937 ( .A(n668), .Y(n667) );
  OAI2B2X1 U3938 ( .A1N(Output2[105]), .A0(n3432), .B0(n3508), .B1(n3433), .Y(
        n668) );
  CLKINVX1 U3939 ( .A(Input2[105]), .Y(n3508) );
  XOR2X1 U3940 ( .A(n3509), .B(n1107), .Y(Output2[105]) );
  CLKINVX1 U3941 ( .A(n3510), .Y(n1107) );
  OAI221X1 U3942 ( .A0(n3511), .A1(n2273), .B0(n2161), .B1(n2274), .C0(n3512), 
        .Y(n3510) );
  AOI2BB2X1 U3943 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[107]), .B1(n294), 
        .A0N(n285), .A1N(n2171), .Y(n3512) );
  XNOR2X1 U3944 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_27_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[107]), .Y(n2171) );
  MXI2X1 U3945 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[111]), .B(n3513), .S0(
        n307), .Y(n2161) );
  XOR2X1 U3946 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[79]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_63_), .Y(n3513) );
  XOR2X1 U3947 ( .A(n2384), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[7]), .Y(
        n3511) );
  XOR2X1 U3948 ( .A(n2215), .B(n2585), .Y(n2384) );
  XOR2X1 U3949 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_57_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[111]), .Y(n2585) );
  CLKINVX1 U3950 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[63]), .Y(n2215) );
  CLKNAND2X2 U3951 ( .A(Input2[105]), .B(n2288), .Y(n3509) );
  OAI221X1 U3952 ( .A0(n671), .A1(n173), .B0(n3514), .B1(n146), .C0(n3515), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_104_N3) );
  AOI22XL U3953 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_104_), 
        .B0(n228), .B1(Input2[104]), .Y(n3515) );
  CLKINVX1 U3954 ( .A(n1109), .Y(n3514) );
  CLKINVX1 U3955 ( .A(n672), .Y(n671) );
  OAI2B2X1 U3956 ( .A1N(Output2[104]), .A0(n3432), .B0(n3516), .B1(n3433), .Y(
        n672) );
  XOR2X1 U3957 ( .A(n1109), .B(n3517), .Y(Output2[104]) );
  NOR2X1 U3958 ( .A(n249), .B(n3516), .Y(n3517) );
  CLKINVX1 U3959 ( .A(Input2[104]), .Y(n3516) );
  OAI221X1 U3960 ( .A0(n2050), .A1(n2274), .B0(n278), .B1(n3518), .C0(n3519), 
        .Y(n1109) );
  AOI22XL U3961 ( .A0(n263), .A1(n3520), .B0(n295), .B1(n3437), .Y(n3519) );
  XNOR2X1 U3962 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_26_), .B(n3518), .Y(
        n3437) );
  XOR2X1 U3963 ( .A(n2503), .B(n2632), .Y(n3520) );
  XOR2X1 U3964 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_0_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[2]), .Y(n2632) );
  XOR2X1 U3965 ( .A(n2593), .B(n2974), .Y(n2503) );
  CLKINVX1 U3966 ( .A(n2095), .Y(n2974) );
  XNOR2X1 U3967 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_14_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[58]), .Y(n2095) );
  XOR2X1 U3968 ( .A(n3474), .B(n2052), .Y(n2593) );
  XOR2X1 U3969 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_26_), .B(n3487), .Y(
        n2052) );
  CLKINVX1 U3970 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[106]), .Y(n3487) );
  CLKINVX1 U3971 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[104]), .Y(n3518) );
  MXI2X1 U3972 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[105]), .B(n3521), .S0(
        n308), .Y(n2050) );
  XOR2X1 U3973 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[73]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_57_), .Y(n3521) );
  OAI221X1 U3974 ( .A0(n3522), .A1(n2300), .B0(n3523), .B1(n2302), .C0(n3524), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_103_N3) );
  AOI22XL U3975 ( .A0(n186), .A1(n675), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1111), .Y(n3524) );
  OAI2B2X1 U3976 ( .A1N(Output2[103]), .A0(n2250), .B0(n3523), .B1(n2252), .Y(
        n675) );
  XOR2X1 U3977 ( .A(n1111), .B(n3525), .Y(Output2[103]) );
  NOR2X1 U3978 ( .A(n249), .B(n3523), .Y(n3525) );
  OAI221X1 U3979 ( .A0(n2060), .A1(n277), .B0(n2267), .B1(n3096), .C0(n3526), 
        .Y(n1111) );
  AOI222XL U3980 ( .A0(n2312), .A1(n2296), .B0(n2258), .B1(n3527), .C0(n264), 
        .C1(n3528), .Y(n3526) );
  XNOR2X1 U3981 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[7]), .B(n2629), .Y(
        n3528) );
  XOR2X1 U3982 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[39]), .B(n2603), .Y(
        n2629) );
  XNOR2X1 U3983 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_23_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[96]), .Y(n2603) );
  XOR2X1 U3984 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[64]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_21_), .Y(n3527) );
  XOR2X1 U3985 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_24_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[96]), .Y(n2296) );
  CLKINVX1 U3986 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[97]), .Y(n3096) );
  CLKINVX1 U3987 ( .A(Input2[103]), .Y(n3523) );
  CLKINVX1 U3988 ( .A(Inst_forkAE_MainPart2_Tag_Reg_Output_103_), .Y(n3522) );
  OAI221X1 U3989 ( .A0(n678), .A1(n173), .B0(n1112), .B1(n146), .C0(n3529), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_102_N3) );
  AOI22XL U3990 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_102_), 
        .B0(n228), .B1(Input2[102]), .Y(n3529) );
  CLKINVX1 U3991 ( .A(n679), .Y(n678) );
  OAI2B2X1 U3992 ( .A1N(Output2[102]), .A0(n2250), .B0(n3530), .B1(n2252), .Y(
        n679) );
  CLKINVX1 U3993 ( .A(Input2[102]), .Y(n3530) );
  XOR2X1 U3994 ( .A(n3531), .B(n1112), .Y(Output2[102]) );
  CLKINVX1 U3995 ( .A(n3532), .Y(n1112) );
  OAI221X1 U3996 ( .A0(n3533), .A1(n2273), .B0(n3534), .B1(n2274), .C0(n3535), 
        .Y(n3532) );
  AOI22XL U3997 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D2[98]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[97]), .B1(n292), .Y(n3535) );
  XOR2X1 U3998 ( .A(n3536), .B(n3537), .Y(n3534) );
  MXI2X1 U3999 ( .A(n3086), .B(n3538), .S0(n311), .Y(n3537) );
  XOR2X1 U4000 ( .A(n3539), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[68]), .Y(
        n3538) );
  OR2X1 U4001 ( .A(n2173), .B(n2054), .Y(n3536) );
  MXI2X1 U4002 ( .A(n3540), .B(n3541), .S0(n309), .Y(n2054) );
  XOR2X1 U4003 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[68]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_22_), .Y(n3541) );
  MXI2X1 U4004 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[103]), .B(n3542), .S0(
        n314), .Y(n2173) );
  XOR2X1 U4005 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[71]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_23_), .Y(n3542) );
  XOR2X1 U4006 ( .A(n2751), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[28]), .Y(
        n3533) );
  XNOR2X1 U4007 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[52]), .B(n2615), .Y(
        n2751) );
  XOR2X1 U4008 ( .A(n3543), .B(n3086), .Y(n2615) );
  CLKINVX1 U4009 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[100]), .Y(n3086) );
  CLKNAND2X2 U4010 ( .A(Input2[102]), .B(n2288), .Y(n3531) );
  OAI221X1 U4011 ( .A0(n682), .A1(n173), .B0(n1113), .B1(n146), .C0(n3544), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_101_N3) );
  AOI22XL U4012 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_101_), 
        .B0(n227), .B1(Input2[101]), .Y(n3544) );
  CLKINVX1 U4013 ( .A(n683), .Y(n682) );
  OAI2B2X1 U4014 ( .A1N(Output2[101]), .A0(n2250), .B0(n3545), .B1(n2252), .Y(
        n683) );
  CLKINVX1 U4015 ( .A(Input2[101]), .Y(n3545) );
  XOR2X1 U4016 ( .A(n3546), .B(n1113), .Y(Output2[101]) );
  CLKINVX1 U4017 ( .A(n3547), .Y(n1113) );
  OAI222X1 U4018 ( .A0(n3548), .A1(n2274), .B0(n3549), .B1(n2273), .C0(n2730), 
        .C1(n2175), .Y(n3547) );
  CLKINVX1 U4019 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[103]), .Y(n2175) );
  XOR2X1 U4020 ( .A(n2867), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[24]), .Y(
        n3549) );
  XNOR2X1 U4021 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[48]), .B(n2639), .Y(
        n2867) );
  XNOR2X1 U4022 ( .A(n3550), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[96]), .Y(
        n2639) );
  XOR2X1 U4023 ( .A(n3551), .B(n3552), .Y(n3548) );
  MXI2X1 U4024 ( .A(n3553), .B(n3554), .S0(n315), .Y(n3552) );
  XOR2X1 U4025 ( .A(n3555), .B(Inst_forkAE_CipherInst_RF_S_MID_D2[64]), .Y(
        n3554) );
  CLKINVX1 U4026 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[96]), .Y(n3553) );
  OR2X1 U4027 ( .A(n2177), .B(n2058), .Y(n3551) );
  MXI2X1 U4028 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[97]), .B(n3556), .S0(
        n316), .Y(n2058) );
  XOR2X1 U4029 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[65]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_17_), .Y(n3556) );
  CLKNAND2X2 U4030 ( .A(Input2[101]), .B(n2288), .Y(n3546) );
  OAI221X1 U4031 ( .A0(n686), .A1(n173), .B0(n3557), .B1(n145), .C0(n3558), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_100_N3) );
  AOI22XL U4032 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_100_), 
        .B0(n227), .B1(Input2[100]), .Y(n3558) );
  CLKINVX1 U4033 ( .A(n1115), .Y(n3557) );
  CLKINVX1 U4034 ( .A(n687), .Y(n686) );
  OAI2B2X1 U4035 ( .A1N(Output2[100]), .A0(n2250), .B0(n3559), .B1(n2252), .Y(
        n687) );
  XOR2X1 U4036 ( .A(n1115), .B(n3560), .Y(Output2[100]) );
  NOR2X1 U4037 ( .A(n249), .B(n3559), .Y(n3560) );
  CLKINVX1 U4038 ( .A(Input2[100]), .Y(n3559) );
  OAI221X1 U4039 ( .A0(n2177), .A1(n2274), .B0(n283), .B1(n2056), .C0(n3561), 
        .Y(n1115) );
  AOI22XL U4040 ( .A0(n263), .A1(n3562), .B0(n295), .B1(n3540), .Y(n3561) );
  XOR2X1 U4041 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_25_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C2[100]), .Y(n3540) );
  XNOR2X1 U4042 ( .A(n2979), .B(n2123), .Y(n3562) );
  XNOR2X1 U4043 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_7_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[27]), .Y(n2123) );
  XNOR2X1 U4044 ( .A(n2654), .B(n2225), .Y(n2979) );
  XNOR2X1 U4045 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_13_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[51]), .Y(n2225) );
  XOR2X1 U4046 ( .A(n3539), .B(n2179), .Y(n2654) );
  XNOR2X1 U4047 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_25_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[99]), .Y(n2179) );
  CLKINVX1 U4048 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[100]), .Y(n2056) );
  MXI2X1 U4049 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[99]), .B(n3563), .S0(
        n306), .Y(n2177) );
  XOR2X1 U4050 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[67]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_19_), .Y(n3563) );
  OAI221X1 U4051 ( .A0(n1035), .A1(n173), .B0(n3564), .B1(n145), .C0(n3565), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_10_N3) );
  AOI22XL U4052 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_10_), 
        .B0(n227), .B1(Input2[10]), .Y(n3565) );
  CLKINVX1 U4053 ( .A(n1267), .Y(n3564) );
  CLKINVX1 U4054 ( .A(n1036), .Y(n1035) );
  OAI2B2X1 U4055 ( .A1N(Output2[10]), .A0(n2379), .B0(n3566), .B1(n2381), .Y(
        n1036) );
  XOR2X1 U4056 ( .A(n1267), .B(n3567), .Y(Output2[10]) );
  NOR2X1 U4057 ( .A(n249), .B(n3566), .Y(n3567) );
  CLKINVX1 U4058 ( .A(Input2[10]), .Y(n3566) );
  OAI221X1 U4059 ( .A0(n2015), .A1(n2274), .B0(n3506), .B1(n2273), .C0(n3568), 
        .Y(n1267) );
  MXI2X1 U4060 ( .A(n3569), .B(n3570), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D2[8]), .Y(n3568) );
  OAI21X1 U4061 ( .A0(n3571), .A1(n281), .B0(n2267), .Y(n3570) );
  NOR2X1 U4062 ( .A(n2139), .B(n2020), .Y(n3571) );
  NOR3X1 U4063 ( .A(n274), .B(n2139), .C(n2020), .Y(n3569) );
  XNOR2X1 U4064 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_2_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[10]), .Y(n2020) );
  CLKINVX1 U4065 ( .A(n2386), .Y(n2139) );
  XOR2X1 U4066 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_3_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[11]), .Y(n2386) );
  XOR2X1 U4067 ( .A(n2092), .B(n2572), .Y(n3506) );
  XNOR2X1 U4068 ( .A(n3572), .B(Inst_forkAE_CipherInst_RF_S_MID_C2[108]), .Y(
        n2572) );
  CLKINVX1 U4069 ( .A(Inst_forkAE_CipherInst_RF_SHIFT2_OUT[42]), .Y(n2092) );
  MXI2X1 U4070 ( .A(n3343), .B(n3573), .S0(n307), .Y(n2015) );
  XOR2X1 U4071 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C2[116]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[26]), .Y(n3573) );
  XOR2X1 U4072 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_3_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[18]), .Y(n3343) );
  OAI221X1 U4073 ( .A0(n1065), .A1(n173), .B0(n1282), .B1(n145), .C0(n3574), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_1_N3) );
  AOI22XL U4074 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_1_), 
        .B0(n227), .B1(Input2[1]), .Y(n3574) );
  AOI22XL U4075 ( .A0(Input2[1]), .A1(n2627), .B0(n1989), .B1(Output2[1]), .Y(
        n1065) );
  XOR2X1 U4076 ( .A(n3575), .B(n1282), .Y(Output2[1]) );
  CLKINVX1 U4077 ( .A(n3576), .Y(n1282) );
  OAI221X1 U4078 ( .A0(n2141), .A1(n2274), .B0(n2287), .B1(n2273), .C0(n3577), 
        .Y(n3576) );
  AOI2BB2X1 U4079 ( .B0(Inst_forkAE_CipherInst_RF_S_MID_D2[3]), .B1(n294), 
        .A0N(n285), .A1N(n2167), .Y(n3577) );
  XNOR2X1 U4080 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_1_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[3]), .Y(n2167) );
  XOR2X1 U4081 ( .A(n2222), .B(n2688), .Y(n2287) );
  XOR2X1 U4082 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_17_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[103]), .Y(n2688) );
  CLKINVX1 U4083 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[55]), .Y(n2222) );
  MXI2X1 U4084 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[7]), .B(n3578), .S0(
        n308), .Y(n2141) );
  XOR2X1 U4085 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[111]), .Y(n3578) );
  CLKNAND2X2 U4086 ( .A(Input2[1]), .B(n2288), .Y(n3575) );
  OAI221X1 U4087 ( .A0(n1068), .A1(n173), .B0(n1284), .B1(n145), .C0(n3579), 
        .Y(Inst_forkAE_CipherInst_RF_RS2_SFF_0_N3) );
  AOI22XL U4088 ( .A0(n199), .A1(Inst_forkAE_MainPart2_Tag_Reg_Output_0_), 
        .B0(n227), .B1(Input2[0]), .Y(n3579) );
  AOI22XL U4089 ( .A0(Input2[0]), .A1(n2627), .B0(n1989), .B1(Output2[0]), .Y(
        n1068) );
  XOR2X1 U4090 ( .A(n3580), .B(n1284), .Y(Output2[0]) );
  AOI221XL U4091 ( .A0(n2634), .A1(n296), .B0(n2872), .B1(n2293), .C0(n3581), 
        .Y(n1284) );
  AO22X1 U4092 ( .A0(n266), .A1(n2297), .B0(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]), .B1(n292), .Y(n3581) );
  XOR2X1 U4093 ( .A(n2696), .B(n3064), .Y(n2297) );
  CLKINVX1 U4094 ( .A(n2102), .Y(n3064) );
  XNOR2X1 U4095 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_12_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[50]), .Y(n2102) );
  XOR2X1 U4096 ( .A(n3555), .B(n2060), .Y(n2696) );
  XNOR2X1 U4097 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_24_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[98]), .Y(n2060) );
  CLKINVX1 U4098 ( .A(n2046), .Y(n2872) );
  MXI2X1 U4099 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[1]), .B(n3582), .S0(
        n311), .Y(n2046) );
  XOR2X1 U4100 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D2[9]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D2[105]), .Y(n3582) );
  XOR2X1 U4101 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX2_0_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT2_OUT[15]), .Y(n2634) );
  CLKNAND2X2 U4102 ( .A(Input2[0]), .B(n2288), .Y(n3580) );
  OAI221X1 U4103 ( .A0(n1389), .A1(n173), .B0(n3583), .B1(n149), .C0(n3584), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_99_N3) );
  AOI22XL U4104 ( .A0(n199), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_99_), 
        .B0(n227), .B1(Input1[99]), .Y(n3584) );
  CLKINVX1 U4105 ( .A(n1810), .Y(n3583) );
  CLKINVX1 U4106 ( .A(n1390), .Y(n1389) );
  OAI2B2X1 U4107 ( .A1N(Output1[99]), .A0(n2250), .B0(n3585), .B1(n2252), .Y(
        n1390) );
  XOR2X1 U4108 ( .A(n1810), .B(n3586), .Y(Output1[99]) );
  NOR2X1 U4109 ( .A(n249), .B(n3585), .Y(n3586) );
  CLKINVX1 U4110 ( .A(Input1[99]), .Y(n3585) );
  OAI2B11X1 U4111 ( .A1N(Inst_forkAE_CipherInst_RF_S_MID_D1[98]), .A0(n2255), 
        .B0(n3587), .C0(n3588), .Y(n1810) );
  AOI22XL U4112 ( .A0(n2258), .A1(n3589), .B0(n261), .B1(n3590), .Y(n3588) );
  XOR2X1 U4113 ( .A(n3591), .B(n3592), .Y(n3590) );
  XOR2X1 U4114 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[66]), .B(n3593), .Y(
        n3589) );
  MXI2X1 U4115 ( .A(n3594), .B(n3595), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[100]), .Y(n3587) );
  OAI21X1 U4116 ( .A0(n3596), .A1(n282), .B0(n2267), .Y(n3595) );
  NOR2X1 U4117 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .Y(n3596) );
  NOR3X1 U4118 ( .A(n274), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .Y(n3594) );
  OAI221X1 U4119 ( .A0(n1393), .A1(n173), .B0(n3597), .B1(n158), .C0(n3598), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_98_N3) );
  AOI22XL U4120 ( .A0(n199), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_98_), 
        .B0(n227), .B1(Input1[98]), .Y(n3598) );
  CLKINVX1 U4121 ( .A(n1812), .Y(n3597) );
  CLKINVX1 U4122 ( .A(n1394), .Y(n1393) );
  OAI2B2X1 U4123 ( .A1N(Output1[98]), .A0(n2250), .B0(n3599), .B1(n2252), .Y(
        n1394) );
  XOR2X1 U4124 ( .A(n1812), .B(n3600), .Y(Output1[98]) );
  NOR2X1 U4125 ( .A(n249), .B(n3599), .Y(n3600) );
  CLKINVX1 U4126 ( .A(Input1[98]), .Y(n3599) );
  OAI221X1 U4127 ( .A0(n3601), .A1(n2273), .B0(n2176), .B1(n2274), .C0(n3602), 
        .Y(n1812) );
  MXI2X1 U4128 ( .A(n3603), .B(n3604), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[96]), .Y(n3602) );
  OAI21X1 U4129 ( .A0(n3605), .A1(n281), .B0(n2267), .Y(n3604) );
  NOR2X1 U4130 ( .A(n2180), .B(n2061), .Y(n3605) );
  NOR3X1 U4131 ( .A(n274), .B(n2180), .C(n2061), .Y(n3603) );
  CLKINVX1 U4132 ( .A(n3606), .Y(n2180) );
  XOR2X1 U4133 ( .A(n3607), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .Y(
        n3601) );
  OAI221X1 U4134 ( .A0(n1397), .A1(n173), .B0(n1813), .B1(n159), .C0(n3608), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_97_N3) );
  AOI22XL U4135 ( .A0(n199), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_97_), 
        .B0(n227), .B1(Input1[97]), .Y(n3608) );
  CLKINVX1 U4136 ( .A(n1398), .Y(n1397) );
  OAI2B2X1 U4137 ( .A1N(Output1[97]), .A0(n2250), .B0(n3609), .B1(n2252), .Y(
        n1398) );
  CLKINVX1 U4138 ( .A(Input1[97]), .Y(n3609) );
  XOR2X1 U4139 ( .A(n3610), .B(n1813), .Y(Output1[97]) );
  CLKINVX1 U4140 ( .A(n3611), .Y(n1813) );
  OAI221X1 U4141 ( .A0(n3612), .A1(n2273), .B0(n2057), .B1(n2274), .C0(n3613), 
        .Y(n3611) );
  AOI22XL U4142 ( .A0(n291), .A1(n2061), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[99]), .B1(n299), .Y(n3613) );
  XOR2X1 U4143 ( .A(n3614), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .Y(
        n3612) );
  CLKNAND2X2 U4144 ( .A(Input1[97]), .B(n2288), .Y(n3610) );
  OAI221X1 U4145 ( .A0(n1401), .A1(n173), .B0(n1814), .B1(n159), .C0(n3615), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_96_N3) );
  AOI22XL U4146 ( .A0(n199), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_96_), 
        .B0(n227), .B1(Input1[96]), .Y(n3615) );
  CLKINVX1 U4147 ( .A(n1402), .Y(n1401) );
  OAI2B2X1 U4148 ( .A1N(Output1[96]), .A0(n2250), .B0(n3616), .B1(n2252), .Y(
        n1402) );
  XNOR2X1 U4149 ( .A(n1814), .B(n3617), .Y(Output1[96]) );
  NOR2X1 U4150 ( .A(n249), .B(n3616), .Y(n3617) );
  CLKINVX1 U4151 ( .A(Input1[96]), .Y(n3616) );
  AOI221XL U4152 ( .A0(n2178), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[96]), .C0(n3618), .Y(n1814) );
  AO22X1 U4153 ( .A0(n266), .A1(n3619), .B0(n300), .B1(n3620), .Y(n3618) );
  XOR2X1 U4154 ( .A(n3621), .B(n2124), .Y(n3619) );
  CLKINVX1 U4155 ( .A(n3622), .Y(n2178) );
  OAI221X1 U4156 ( .A0(n3623), .A1(n2300), .B0(n3624), .B1(n2302), .C0(n3625), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_95_N3) );
  AOI22XL U4157 ( .A0(n186), .A1(n1405), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1816), .Y(n3625) );
  OAI222X1 U4158 ( .A0(n2304), .A1(n3626), .B0(n3627), .B1(n3628), .C0(n3624), 
        .C1(n2305), .Y(n1405) );
  CLKINVX1 U4159 ( .A(Output1[95]), .Y(n3626) );
  XOR2X1 U4160 ( .A(n1816), .B(n3629), .Y(Output1[95]) );
  NOR2X1 U4161 ( .A(n249), .B(n3624), .Y(n3629) );
  OAI221X1 U4162 ( .A0(n3630), .A1(n2273), .B0(n2267), .B1(n3631), .C0(n3632), 
        .Y(n1816) );
  AOI222XL U4163 ( .A0(n291), .A1(n2188), .B0(n2258), .B1(n3633), .C0(n2312), 
        .C1(n3634), .Y(n3632) );
  XOR2X1 U4164 ( .A(n3635), .B(n3636), .Y(n3633) );
  XOR2X1 U4165 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[48]), .B(n3637), .Y(
        n3636) );
  CLKINVX1 U4166 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .Y(n3631) );
  CLKINVX1 U4167 ( .A(Input1[95]), .Y(n3624) );
  CLKINVX1 U4168 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_95_), .Y(n3623) );
  OAI221X1 U4169 ( .A0(n1408), .A1(n172), .B0(n1817), .B1(n159), .C0(n3638), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_94_N3) );
  AOI22XL U4170 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_94_), 
        .B0(n227), .B1(Input1[94]), .Y(n3638) );
  CLKINVX1 U4171 ( .A(n1409), .Y(n1408) );
  OAI2B2X1 U4172 ( .A1N(Output1[94]), .A0(n2304), .B0(n3639), .B1(n2305), .Y(
        n1409) );
  CLKINVX1 U4173 ( .A(Input1[94]), .Y(n3639) );
  XOR2X1 U4174 ( .A(n3640), .B(n1817), .Y(Output1[94]) );
  CLKINVX1 U4175 ( .A(n3641), .Y(n1817) );
  OAI221X1 U4176 ( .A0(n3642), .A1(n2274), .B0(n3643), .B1(n2273), .C0(n3644), 
        .Y(n3641) );
  AOI22XL U4177 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[90]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .B1(n291), .Y(n3644) );
  XOR2X1 U4178 ( .A(n3645), .B(n3646), .Y(n3642) );
  MXI2X1 U4179 ( .A(n3647), .B(n3648), .S0(n309), .Y(n3646) );
  XOR2X1 U4180 ( .A(n3649), .B(n3650), .Y(n3648) );
  XOR2X1 U4181 ( .A(n3651), .B(n3652), .Y(n3649) );
  CLKNAND2X2 U4182 ( .A(n2184), .B(n3653), .Y(n3645) );
  CLKNAND2X2 U4183 ( .A(Input1[94]), .B(n2288), .Y(n3640) );
  OAI221X1 U4184 ( .A0(n1412), .A1(n172), .B0(n3654), .B1(n159), .C0(n3655), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_93_N3) );
  AOI22XL U4185 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_93_), 
        .B0(n227), .B1(Input1[93]), .Y(n3655) );
  CLKINVX1 U4186 ( .A(n1819), .Y(n3654) );
  CLKINVX1 U4187 ( .A(n1413), .Y(n1412) );
  OAI2B2X1 U4188 ( .A1N(Output1[93]), .A0(n2304), .B0(n3656), .B1(n2305), .Y(
        n1413) );
  XOR2X1 U4189 ( .A(n1819), .B(n3657), .Y(Output1[93]) );
  NOR2X1 U4190 ( .A(n249), .B(n3656), .Y(n3657) );
  CLKINVX1 U4191 ( .A(Input1[93]), .Y(n3656) );
  OAI222X1 U4192 ( .A0(n2730), .A1(n3658), .B0(n3659), .B1(n2274), .C0(n3660), 
        .C1(n2273), .Y(n1819) );
  XOR2X1 U4193 ( .A(n3661), .B(n3662), .Y(n3659) );
  MXI2X1 U4194 ( .A(n3663), .B(n3664), .S0(n310), .Y(n3662) );
  XOR2X1 U4195 ( .A(n3665), .B(n3666), .Y(n3664) );
  XOR2X1 U4196 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .B(n3667), .Y(
        n3666) );
  XOR2X1 U4197 ( .A(n1991), .B(n3668), .Y(n3665) );
  CLKNAND2X2 U4198 ( .A(n3669), .B(n3670), .Y(n3661) );
  CLKINVX1 U4199 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .Y(n3658) );
  OAI221X1 U4200 ( .A0(n1416), .A1(n172), .B0(n1821), .B1(n159), .C0(n3671), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_92_N3) );
  AOI22XL U4201 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_92_), 
        .B0(n227), .B1(Input1[92]), .Y(n3671) );
  CLKINVX1 U4202 ( .A(n1417), .Y(n1416) );
  OAI2B2X1 U4203 ( .A1N(Input1[92]), .A0(n2305), .B0(n3672), .B1(n2304), .Y(
        n1417) );
  CLKINVX1 U4204 ( .A(Output1[92]), .Y(n3672) );
  XOR2X1 U4205 ( .A(n3673), .B(n1821), .Y(Output1[92]) );
  AOI221XL U4206 ( .A0(n3674), .A1(n296), .B0(n2066), .B1(n2293), .C0(n3675), 
        .Y(n1821) );
  AO22X1 U4207 ( .A0(n266), .A1(n3676), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .B1(n292), .Y(n3675) );
  CLKINVX1 U4208 ( .A(n3669), .Y(n2066) );
  MXI2X1 U4209 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[91]), .B(n3677), .S0(
        n314), .Y(n3669) );
  XOR2X1 U4210 ( .A(n3678), .B(n3679), .Y(n3677) );
  XOR2X1 U4211 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[51]), .B(n3680), .Y(
        n3679) );
  CLKNAND2X2 U4212 ( .A(Input1[92]), .B(n2288), .Y(n3673) );
  OAI221X1 U4213 ( .A0(n1420), .A1(n172), .B0(n3681), .B1(n159), .C0(n3682), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_91_N3) );
  AOI22XL U4214 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_91_), 
        .B0(n227), .B1(Input1[91]), .Y(n3682) );
  CLKINVX1 U4215 ( .A(n1823), .Y(n3681) );
  CLKINVX1 U4216 ( .A(n1421), .Y(n1420) );
  OAI2B2X1 U4217 ( .A1N(Output1[91]), .A0(n2304), .B0(n3683), .B1(n2305), .Y(
        n1421) );
  XOR2X1 U4218 ( .A(n1823), .B(n3684), .Y(Output1[91]) );
  NOR2X1 U4219 ( .A(n250), .B(n3683), .Y(n3684) );
  CLKINVX1 U4220 ( .A(Input1[91]), .Y(n3683) );
  OAI211XL U4221 ( .A0(n3685), .A1(n2273), .B0(n3686), .C0(n3687), .Y(n1823)
         );
  AOI22XL U4222 ( .A0(n2258), .A1(n3688), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[90]), .B1(n2312), .Y(n3687) );
  XNOR2X1 U4223 ( .A(n3689), .B(n3690), .Y(n3688) );
  XOR2X1 U4224 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[50]), .B(n3691), .Y(
        n3690) );
  MXI2X1 U4225 ( .A(n3692), .B(n3693), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[92]), .Y(n3686) );
  OAI21X1 U4226 ( .A0(n3694), .A1(n281), .B0(n2267), .Y(n3693) );
  NOR2X1 U4227 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .Y(n3694) );
  NOR3X1 U4228 ( .A(n274), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .Y(n3692) );
  OAI221X1 U4229 ( .A0(n1424), .A1(n172), .B0(n3695), .B1(n159), .C0(n3696), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_90_N3) );
  AOI22XL U4230 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_90_), 
        .B0(n226), .B1(Input1[90]), .Y(n3696) );
  CLKINVX1 U4231 ( .A(n1825), .Y(n3695) );
  CLKINVX1 U4232 ( .A(n1425), .Y(n1424) );
  OAI2B2X1 U4233 ( .A1N(Output1[90]), .A0(n2304), .B0(n3697), .B1(n2305), .Y(
        n1425) );
  XOR2X1 U4234 ( .A(n1825), .B(n3698), .Y(Output1[90]) );
  NOR2X1 U4235 ( .A(n250), .B(n3697), .Y(n3698) );
  CLKINVX1 U4236 ( .A(Input1[90]), .Y(n3697) );
  OAI221X1 U4237 ( .A0(n2184), .A1(n2274), .B0(n3699), .B1(n2273), .C0(n3700), 
        .Y(n1825) );
  MXI2X1 U4238 ( .A(n3701), .B(n3702), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[88]), .Y(n3700) );
  OAI21X1 U4239 ( .A0(n3703), .A1(n282), .B0(n2267), .Y(n3702) );
  NOR2X1 U4240 ( .A(n2068), .B(n2188), .Y(n3703) );
  NOR3X1 U4241 ( .A(n275), .B(n2188), .C(n2068), .Y(n3701) );
  MXI2X1 U4242 ( .A(n3674), .B(n3704), .S0(n315), .Y(n2184) );
  XOR2X1 U4243 ( .A(n3705), .B(n3706), .Y(n3704) );
  XOR2X1 U4244 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .B(n3707), .Y(
        n3706) );
  XOR2X1 U4245 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_23_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .Y(n3674) );
  OAI221X1 U4246 ( .A0(n1738), .A1(n172), .B0(n1954), .B1(n159), .C0(n3708), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_9_N3) );
  AOI22XL U4247 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_9_), 
        .B0(n226), .B1(Input1[9]), .Y(n3708) );
  CLKINVX1 U4248 ( .A(n1739), .Y(n1738) );
  OAI2B2X1 U4249 ( .A1N(Input1[9]), .A0(n2381), .B0(n3709), .B1(n2379), .Y(
        n1739) );
  CLKINVX1 U4250 ( .A(Output1[9]), .Y(n3709) );
  XOR2X1 U4251 ( .A(n3710), .B(n1954), .Y(Output1[9]) );
  AOI221XL U4252 ( .A0(n2016), .A1(n2293), .B0(n261), .B1(n3711), .C0(n3712), 
        .Y(n1954) );
  AO22X1 U4253 ( .A0(n292), .A1(n2021), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[11]), .B1(n301), .Y(n3712) );
  CLKINVX1 U4254 ( .A(n3713), .Y(n2016) );
  CLKNAND2X2 U4255 ( .A(Input1[9]), .B(n2288), .Y(n3710) );
  OAI221X1 U4256 ( .A0(n1428), .A1(n172), .B0(n1826), .B1(n159), .C0(n3714), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_89_N3) );
  AOI22XL U4257 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_89_), 
        .B0(n226), .B1(Input1[89]), .Y(n3714) );
  CLKINVX1 U4258 ( .A(n1429), .Y(n1428) );
  OAI2B2X1 U4259 ( .A1N(Output1[89]), .A0(n2304), .B0(n3715), .B1(n2305), .Y(
        n1429) );
  XNOR2X1 U4260 ( .A(n1826), .B(n3716), .Y(Output1[89]) );
  NOR2X1 U4261 ( .A(n250), .B(n3715), .Y(n3716) );
  CLKINVX1 U4262 ( .A(Input1[89]), .Y(n3715) );
  AOI221XL U4263 ( .A0(n2063), .A1(n2293), .B0(n2068), .B1(n291), .C0(n3717), 
        .Y(n1826) );
  AO22X1 U4264 ( .A0(n3718), .A1(n268), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[91]), .B1(n301), .Y(n3717) );
  CLKINVX1 U4265 ( .A(n3653), .Y(n2063) );
  MXI2X1 U4266 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .B(n3719), .S0(
        n316), .Y(n3653) );
  XOR2X1 U4267 ( .A(n3720), .B(n3721), .Y(n3719) );
  XOR2X1 U4268 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .B(n3722), .Y(
        n3721) );
  OAI221X1 U4269 ( .A0(n1432), .A1(n172), .B0(n1828), .B1(n159), .C0(n3723), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_88_N3) );
  AOI22XL U4270 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_88_), 
        .B0(n226), .B1(Input1[88]), .Y(n3723) );
  CLKINVX1 U4271 ( .A(n1433), .Y(n1432) );
  OAI2B2X1 U4272 ( .A1N(Input1[88]), .A0(n2305), .B0(n3724), .B1(n2304), .Y(
        n1433) );
  CLKNAND2X2 U4273 ( .A(dec), .B(n3627), .Y(n2304) );
  CLKINVX1 U4274 ( .A(Output1[88]), .Y(n3724) );
  XOR2X1 U4275 ( .A(n3725), .B(n1828), .Y(Output1[88]) );
  AOI221XL U4276 ( .A0(n3634), .A1(n297), .B0(n2186), .B1(n2293), .C0(n3726), 
        .Y(n1828) );
  AO22X1 U4277 ( .A0(n266), .A1(n3727), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[88]), .B1(n292), .Y(n3726) );
  CLKINVX1 U4278 ( .A(n3670), .Y(n2186) );
  MXI2X1 U4279 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .B(n3728), .S0(
        n313), .Y(n3670) );
  XOR2X1 U4280 ( .A(n3729), .B(n3730), .Y(n3728) );
  XOR2X1 U4281 ( .A(n1992), .B(n3731), .Y(n3730) );
  XOR2X1 U4282 ( .A(n3732), .B(n3733), .Y(n3729) );
  XOR2X1 U4283 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_22_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[88]), .Y(n3634) );
  CLKNAND2X2 U4284 ( .A(Input1[88]), .B(n2288), .Y(n3725) );
  CLKNAND2X2 U4285 ( .A(n3627), .B(n3734), .Y(n2305) );
  OAI221X1 U4286 ( .A0(n3735), .A1(n2300), .B0(n3736), .B1(n2302), .C0(n3737), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_87_N3) );
  AOI22XL U4287 ( .A0(n186), .A1(n1436), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1830), .Y(n3737) );
  OAI222X1 U4288 ( .A0(n2407), .A1(n3738), .B0(n3739), .B1(n3740), .C0(n3736), 
        .C1(n2408), .Y(n1436) );
  CLKINVX1 U4289 ( .A(Output1[87]), .Y(n3738) );
  XOR2X1 U4290 ( .A(n1830), .B(n3741), .Y(Output1[87]) );
  NOR2X1 U4291 ( .A(n250), .B(n3736), .Y(n3741) );
  OAI221X1 U4292 ( .A0(n3742), .A1(n2273), .B0(n2267), .B1(n3743), .C0(n3744), 
        .Y(n1830) );
  AOI222XL U4293 ( .A0(n291), .A1(n2196), .B0(n2258), .B1(n3745), .C0(n2312), 
        .C1(n3746), .Y(n3744) );
  XOR2X1 U4294 ( .A(n3747), .B(n3748), .Y(n3745) );
  XOR2X1 U4295 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[40]), .B(n3749), .Y(
        n3748) );
  CLKINVX1 U4296 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .Y(n3743) );
  CLKINVX1 U4297 ( .A(Input1[87]), .Y(n3736) );
  CLKINVX1 U4298 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_87_), .Y(n3735) );
  OAI221X1 U4299 ( .A0(n1439), .A1(n172), .B0(n1831), .B1(n158), .C0(n3750), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_86_N3) );
  AOI22XL U4300 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_86_), 
        .B0(n226), .B1(Input1[86]), .Y(n3750) );
  CLKINVX1 U4301 ( .A(n1440), .Y(n1439) );
  OAI2B2X1 U4302 ( .A1N(Output1[86]), .A0(n2407), .B0(n3751), .B1(n2408), .Y(
        n1440) );
  CLKINVX1 U4303 ( .A(Input1[86]), .Y(n3751) );
  XOR2X1 U4304 ( .A(n3752), .B(n1831), .Y(Output1[86]) );
  CLKINVX1 U4305 ( .A(n3753), .Y(n1831) );
  OAI221X1 U4306 ( .A0(n3754), .A1(n2274), .B0(n3755), .B1(n2273), .C0(n3756), 
        .Y(n3753) );
  AOI22XL U4307 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[82]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .B1(n291), .Y(n3756) );
  XOR2X1 U4308 ( .A(n3757), .B(n3758), .Y(n3754) );
  MXI2X1 U4309 ( .A(n3759), .B(n3760), .S0(n312), .Y(n3758) );
  XOR2X1 U4310 ( .A(n3761), .B(n3762), .Y(n3760) );
  XNOR2X1 U4311 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .B(n3763), .Y(
        n3761) );
  CLKNAND2X2 U4312 ( .A(n2192), .B(n3764), .Y(n3757) );
  CLKNAND2X2 U4313 ( .A(Input1[86]), .B(n2288), .Y(n3752) );
  OAI221X1 U4314 ( .A0(n1443), .A1(n172), .B0(n3765), .B1(n159), .C0(n3766), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_85_N3) );
  AOI22XL U4315 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_85_), 
        .B0(n226), .B1(Input1[85]), .Y(n3766) );
  CLKINVX1 U4316 ( .A(n1833), .Y(n3765) );
  CLKINVX1 U4317 ( .A(n1444), .Y(n1443) );
  OAI2B2X1 U4318 ( .A1N(Output1[85]), .A0(n2407), .B0(n3767), .B1(n2408), .Y(
        n1444) );
  XOR2X1 U4319 ( .A(n1833), .B(n3768), .Y(Output1[85]) );
  NOR2X1 U4320 ( .A(n250), .B(n3767), .Y(n3768) );
  CLKINVX1 U4321 ( .A(Input1[85]), .Y(n3767) );
  OAI222X1 U4322 ( .A0(n2730), .A1(n3769), .B0(n3770), .B1(n2274), .C0(n3771), 
        .C1(n2273), .Y(n1833) );
  XOR2X1 U4323 ( .A(n3772), .B(n3773), .Y(n3770) );
  MXI2X1 U4324 ( .A(n3774), .B(n3775), .S0(n313), .Y(n3773) );
  XOR2X1 U4325 ( .A(n3776), .B(n3777), .Y(n3775) );
  XNOR2X1 U4326 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .B(n3778), .Y(
        n3776) );
  CLKNAND2X2 U4327 ( .A(n3779), .B(n3780), .Y(n3772) );
  CLKINVX1 U4328 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .Y(n3769) );
  OAI221X1 U4329 ( .A0(n1447), .A1(n172), .B0(n1835), .B1(n158), .C0(n3781), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_84_N3) );
  AOI22XL U4330 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_84_), 
        .B0(n226), .B1(Input1[84]), .Y(n3781) );
  CLKINVX1 U4331 ( .A(n1448), .Y(n1447) );
  OAI2B2X1 U4332 ( .A1N(Input1[84]), .A0(n2408), .B0(n3782), .B1(n2407), .Y(
        n1448) );
  CLKINVX1 U4333 ( .A(Output1[84]), .Y(n3782) );
  XOR2X1 U4334 ( .A(n3783), .B(n1835), .Y(Output1[84]) );
  AOI221XL U4335 ( .A0(n3784), .A1(n297), .B0(n2073), .B1(n2293), .C0(n3785), 
        .Y(n1835) );
  AO22X1 U4336 ( .A0(n267), .A1(n3786), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .B1(n292), .Y(n3785) );
  CLKINVX1 U4337 ( .A(n3779), .Y(n2073) );
  MXI2X1 U4338 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[83]), .B(n3787), .S0(
        n312), .Y(n3779) );
  XOR2X1 U4339 ( .A(n3788), .B(n3789), .Y(n3787) );
  XOR2X1 U4340 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[43]), .B(n3790), .Y(
        n3789) );
  CLKNAND2X2 U4341 ( .A(Input1[84]), .B(n2288), .Y(n3783) );
  OAI221X1 U4342 ( .A0(n1451), .A1(n172), .B0(n3791), .B1(n158), .C0(n3792), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_83_N3) );
  AOI22XL U4343 ( .A0(n198), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_83_), 
        .B0(n226), .B1(Input1[83]), .Y(n3792) );
  CLKINVX1 U4344 ( .A(n1837), .Y(n3791) );
  CLKINVX1 U4345 ( .A(n1452), .Y(n1451) );
  OAI2B2X1 U4346 ( .A1N(Output1[83]), .A0(n2407), .B0(n3793), .B1(n2408), .Y(
        n1452) );
  XOR2X1 U4347 ( .A(n1837), .B(n3794), .Y(Output1[83]) );
  NOR2X1 U4348 ( .A(n250), .B(n3793), .Y(n3794) );
  CLKINVX1 U4349 ( .A(Input1[83]), .Y(n3793) );
  OAI211XL U4350 ( .A0(n3795), .A1(n2273), .B0(n3796), .C0(n3797), .Y(n1837)
         );
  AOI22XL U4351 ( .A0(n2258), .A1(n3798), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[82]), .B1(n2312), .Y(n3797) );
  XNOR2X1 U4352 ( .A(n3799), .B(n3800), .Y(n3798) );
  XOR2X1 U4353 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[42]), .B(n3801), .Y(
        n3800) );
  MXI2X1 U4354 ( .A(n3802), .B(n3803), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[84]), .Y(n3796) );
  OAI21X1 U4355 ( .A0(n3804), .A1(n281), .B0(n2267), .Y(n3803) );
  NOR2X1 U4356 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .Y(n3804) );
  NOR3X1 U4357 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .Y(n3802) );
  OAI221X1 U4358 ( .A0(n1455), .A1(n171), .B0(n3805), .B1(n158), .C0(n3806), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_82_N3) );
  AOI22XL U4359 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_82_), 
        .B0(n226), .B1(Input1[82]), .Y(n3806) );
  CLKINVX1 U4360 ( .A(n1839), .Y(n3805) );
  CLKINVX1 U4361 ( .A(n1456), .Y(n1455) );
  OAI2B2X1 U4362 ( .A1N(Output1[82]), .A0(n2407), .B0(n3807), .B1(n2408), .Y(
        n1456) );
  XOR2X1 U4363 ( .A(n1839), .B(n3808), .Y(Output1[82]) );
  NOR2X1 U4364 ( .A(n250), .B(n3807), .Y(n3808) );
  CLKINVX1 U4365 ( .A(Input1[82]), .Y(n3807) );
  OAI221X1 U4366 ( .A0(n2192), .A1(n2274), .B0(n3809), .B1(n2273), .C0(n3810), 
        .Y(n1839) );
  MXI2X1 U4367 ( .A(n3811), .B(n3812), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[80]), .Y(n3810) );
  OAI21X1 U4368 ( .A0(n3813), .A1(n282), .B0(n2267), .Y(n3812) );
  NOR2X1 U4369 ( .A(n2075), .B(n2196), .Y(n3813) );
  NOR3X1 U4370 ( .A(n275), .B(n2196), .C(n2075), .Y(n3811) );
  MXI2X1 U4371 ( .A(n3784), .B(n3814), .S0(n314), .Y(n2192) );
  XOR2X1 U4372 ( .A(n3815), .B(n3816), .Y(n3814) );
  XOR2X1 U4373 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .B(n3817), .Y(
        n3816) );
  XOR2X1 U4374 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_21_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .Y(n3784) );
  OAI221X1 U4375 ( .A0(n1459), .A1(n171), .B0(n1840), .B1(n158), .C0(n3818), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_81_N3) );
  AOI22XL U4376 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_81_), 
        .B0(n226), .B1(Input1[81]), .Y(n3818) );
  CLKINVX1 U4377 ( .A(n1460), .Y(n1459) );
  OAI2B2X1 U4378 ( .A1N(Output1[81]), .A0(n2407), .B0(n3819), .B1(n2408), .Y(
        n1460) );
  XNOR2X1 U4379 ( .A(n1840), .B(n3820), .Y(Output1[81]) );
  NOR2X1 U4380 ( .A(n250), .B(n3819), .Y(n3820) );
  CLKINVX1 U4381 ( .A(Input1[81]), .Y(n3819) );
  AOI221XL U4382 ( .A0(n2070), .A1(n2293), .B0(n2075), .B1(n291), .C0(n3821), 
        .Y(n1840) );
  AO22X1 U4383 ( .A0(n267), .A1(n3822), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[83]), .B1(n302), .Y(n3821) );
  CLKINVX1 U4384 ( .A(n3764), .Y(n2070) );
  MXI2X1 U4385 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .B(n3823), .S0(
        n315), .Y(n3764) );
  XOR2X1 U4386 ( .A(n3824), .B(n3825), .Y(n3823) );
  XOR2X1 U4387 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .B(n3826), .Y(
        n3825) );
  OAI221X1 U4388 ( .A0(n1463), .A1(n171), .B0(n1842), .B1(n158), .C0(n3827), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_80_N3) );
  AOI22XL U4389 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_80_), 
        .B0(n226), .B1(Input1[80]), .Y(n3827) );
  CLKINVX1 U4390 ( .A(n1464), .Y(n1463) );
  OAI2B2X1 U4391 ( .A1N(Input1[80]), .A0(n2408), .B0(n3828), .B1(n2407), .Y(
        n1464) );
  CLKNAND2X2 U4392 ( .A(dec), .B(n3739), .Y(n2407) );
  CLKINVX1 U4393 ( .A(Output1[80]), .Y(n3828) );
  XOR2X1 U4394 ( .A(n3829), .B(n1842), .Y(Output1[80]) );
  AOI221XL U4395 ( .A0(n3746), .A1(n297), .B0(n2194), .B1(n2293), .C0(n3830), 
        .Y(n1842) );
  AO22X1 U4396 ( .A0(n267), .A1(n3831), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[80]), .B1(n292), .Y(n3830) );
  CLKINVX1 U4397 ( .A(n3780), .Y(n2194) );
  MXI2X1 U4398 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .B(n3832), .S0(
        n316), .Y(n3780) );
  XNOR2X1 U4399 ( .A(n3833), .B(n3834), .Y(n3832) );
  XOR2X1 U4400 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[41]), .B(n3835), .Y(
        n3834) );
  XOR2X1 U4401 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_20_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[80]), .Y(n3746) );
  CLKNAND2X2 U4402 ( .A(Input1[80]), .B(n2288), .Y(n3829) );
  CLKNAND2X2 U4403 ( .A(n3739), .B(n3734), .Y(n2408) );
  AO21X1 U4404 ( .A0(Block_Size[2]), .A1(Block_Size[0]), .B0(n3836), .Y(n3739)
         );
  OAI221X1 U4405 ( .A0(n1742), .A1(n171), .B0(n1956), .B1(n158), .C0(n3837), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_8_N3) );
  AOI22XL U4406 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_8_), 
        .B0(n226), .B1(Input1[8]), .Y(n3837) );
  CLKINVX1 U4407 ( .A(n1743), .Y(n1742) );
  OAI2B2X1 U4408 ( .A1N(Input1[8]), .A0(n2381), .B0(n3838), .B1(n2379), .Y(
        n1743) );
  CLKINVX1 U4409 ( .A(Output1[8]), .Y(n3838) );
  XOR2X1 U4410 ( .A(n3839), .B(n1956), .Y(Output1[8]) );
  AOI221XL U4411 ( .A0(n3840), .A1(n297), .B0(n2138), .B1(n2293), .C0(n3841), 
        .Y(n1956) );
  OAI2BB2X1 U4412 ( .B0(n3842), .B1(n284), .A0N(n3843), .A1N(n269), .Y(n3841)
         );
  CLKINVX1 U4413 ( .A(n3844), .Y(n2138) );
  CLKNAND2X2 U4414 ( .A(Input1[8]), .B(n2288), .Y(n3839) );
  OAI221X1 U4415 ( .A0(n3845), .A1(n2300), .B0(n3846), .B1(n2302), .C0(n3847), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_79_N3) );
  AOI22XL U4416 ( .A0(n186), .A1(n1467), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1844), .Y(n3847) );
  OAI222X1 U4417 ( .A0(n2507), .A1(n3848), .B0(n3740), .B1(n3849), .C0(n3846), 
        .C1(n2508), .Y(n1467) );
  CLKINVX1 U4418 ( .A(Output1[79]), .Y(n3848) );
  XOR2X1 U4419 ( .A(n1844), .B(n3850), .Y(Output1[79]) );
  NOR2X1 U4420 ( .A(n250), .B(n3846), .Y(n3850) );
  OAI221X1 U4421 ( .A0(n3851), .A1(n2273), .B0(n2267), .B1(n3852), .C0(n3853), 
        .Y(n1844) );
  AOI222XL U4422 ( .A0(n291), .A1(n2204), .B0(n2258), .B1(n3854), .C0(n2312), 
        .C1(n3855), .Y(n3853) );
  XOR2X1 U4423 ( .A(n3856), .B(n3857), .Y(n3854) );
  XOR2X1 U4424 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[32]), .B(n3858), .Y(
        n3857) );
  CLKINVX1 U4425 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .Y(n3852) );
  CLKINVX1 U4426 ( .A(Input1[79]), .Y(n3846) );
  CLKINVX1 U4427 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_79_), .Y(n3845) );
  OAI221X1 U4428 ( .A0(n1470), .A1(n171), .B0(n1845), .B1(n158), .C0(n3859), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_78_N3) );
  AOI22XL U4429 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_78_), 
        .B0(n226), .B1(Input1[78]), .Y(n3859) );
  CLKINVX1 U4430 ( .A(n1471), .Y(n1470) );
  OAI2B2X1 U4431 ( .A1N(Output1[78]), .A0(n2507), .B0(n3860), .B1(n2508), .Y(
        n1471) );
  CLKINVX1 U4432 ( .A(Input1[78]), .Y(n3860) );
  XOR2X1 U4433 ( .A(n3861), .B(n1845), .Y(Output1[78]) );
  CLKINVX1 U4434 ( .A(n3862), .Y(n1845) );
  OAI221X1 U4435 ( .A0(n3863), .A1(n2274), .B0(n3864), .B1(n2273), .C0(n3865), 
        .Y(n3862) );
  AOI22XL U4436 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[74]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .B1(n291), .Y(n3865) );
  XOR2X1 U4437 ( .A(n3866), .B(n3867), .Y(n3863) );
  MXI2X1 U4438 ( .A(n3868), .B(n3869), .S0(n312), .Y(n3867) );
  XOR2X1 U4439 ( .A(n3870), .B(n3871), .Y(n3869) );
  XNOR2X1 U4440 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .B(n3872), .Y(
        n3870) );
  CLKNAND2X2 U4441 ( .A(n2200), .B(n3873), .Y(n3866) );
  CLKNAND2X2 U4442 ( .A(Input1[78]), .B(n2288), .Y(n3861) );
  OAI221X1 U4443 ( .A0(n1474), .A1(n171), .B0(n3874), .B1(n158), .C0(n3875), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_77_N3) );
  AOI22XL U4444 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_77_), 
        .B0(n225), .B1(Input1[77]), .Y(n3875) );
  CLKINVX1 U4445 ( .A(n1847), .Y(n3874) );
  CLKINVX1 U4446 ( .A(n1475), .Y(n1474) );
  OAI2B2X1 U4447 ( .A1N(Output1[77]), .A0(n2507), .B0(n3876), .B1(n2508), .Y(
        n1475) );
  XOR2X1 U4448 ( .A(n1847), .B(n3877), .Y(Output1[77]) );
  NOR2X1 U4449 ( .A(n250), .B(n3876), .Y(n3877) );
  CLKINVX1 U4450 ( .A(Input1[77]), .Y(n3876) );
  OAI222X1 U4451 ( .A0(n2730), .A1(n3878), .B0(n3879), .B1(n2274), .C0(n3880), 
        .C1(n2273), .Y(n1847) );
  XOR2X1 U4452 ( .A(n3881), .B(n3882), .Y(n3879) );
  MXI2X1 U4453 ( .A(n3883), .B(n3884), .S0(n306), .Y(n3882) );
  XOR2X1 U4454 ( .A(n3885), .B(n3886), .Y(n3884) );
  XNOR2X1 U4455 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .B(n3887), .Y(
        n3885) );
  CLKNAND2X2 U4456 ( .A(n3888), .B(n3889), .Y(n3881) );
  CLKINVX1 U4457 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .Y(n3878) );
  OAI221X1 U4458 ( .A0(n1478), .A1(n171), .B0(n1849), .B1(n158), .C0(n3890), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_76_N3) );
  AOI22XL U4459 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_76_), 
        .B0(n225), .B1(Input1[76]), .Y(n3890) );
  CLKINVX1 U4460 ( .A(n1479), .Y(n1478) );
  OAI2B2X1 U4461 ( .A1N(Input1[76]), .A0(n2508), .B0(n3891), .B1(n2507), .Y(
        n1479) );
  CLKINVX1 U4462 ( .A(Output1[76]), .Y(n3891) );
  XOR2X1 U4463 ( .A(n3892), .B(n1849), .Y(Output1[76]) );
  AOI221XL U4464 ( .A0(n3893), .A1(n297), .B0(n2080), .B1(n2293), .C0(n3894), 
        .Y(n1849) );
  AO22X1 U4465 ( .A0(n267), .A1(n3895), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .B1(n292), .Y(n3894) );
  CLKINVX1 U4466 ( .A(n3888), .Y(n2080) );
  MXI2X1 U4467 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[75]), .B(n3896), .S0(
        n307), .Y(n3888) );
  XOR2X1 U4468 ( .A(n3897), .B(n3898), .Y(n3896) );
  XOR2X1 U4469 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[35]), .B(n3899), .Y(
        n3898) );
  CLKNAND2X2 U4470 ( .A(Input1[76]), .B(n2288), .Y(n3892) );
  OAI221X1 U4471 ( .A0(n1482), .A1(n171), .B0(n3900), .B1(n158), .C0(n3901), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_75_N3) );
  AOI22XL U4472 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_75_), 
        .B0(n225), .B1(Input1[75]), .Y(n3901) );
  CLKINVX1 U4473 ( .A(n1851), .Y(n3900) );
  CLKINVX1 U4474 ( .A(n1483), .Y(n1482) );
  OAI2B2X1 U4475 ( .A1N(Output1[75]), .A0(n2507), .B0(n3902), .B1(n2508), .Y(
        n1483) );
  XOR2X1 U4476 ( .A(n1851), .B(n3903), .Y(Output1[75]) );
  NOR2X1 U4477 ( .A(n250), .B(n3902), .Y(n3903) );
  CLKINVX1 U4478 ( .A(Input1[75]), .Y(n3902) );
  OAI211XL U4479 ( .A0(n3904), .A1(n2273), .B0(n3905), .C0(n3906), .Y(n1851)
         );
  AOI22XL U4480 ( .A0(n2258), .A1(n3907), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[74]), .B1(n2312), .Y(n3906) );
  XNOR2X1 U4481 ( .A(n3908), .B(n3909), .Y(n3907) );
  XOR2X1 U4482 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[34]), .B(n3910), .Y(
        n3909) );
  MXI2X1 U4483 ( .A(n3911), .B(n3912), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[76]), .Y(n3905) );
  OAI21X1 U4484 ( .A0(n3913), .A1(n282), .B0(n2267), .Y(n3912) );
  NOR2X1 U4485 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .Y(n3913) );
  NOR3X1 U4486 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .Y(n3911) );
  OAI221X1 U4487 ( .A0(n1486), .A1(n171), .B0(n3914), .B1(n158), .C0(n3915), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_74_N3) );
  AOI22XL U4488 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_74_), 
        .B0(n225), .B1(Input1[74]), .Y(n3915) );
  CLKINVX1 U4489 ( .A(n1853), .Y(n3914) );
  CLKINVX1 U4490 ( .A(n1487), .Y(n1486) );
  OAI2B2X1 U4491 ( .A1N(Output1[74]), .A0(n2507), .B0(n3916), .B1(n2508), .Y(
        n1487) );
  XOR2X1 U4492 ( .A(n1853), .B(n3917), .Y(Output1[74]) );
  NOR2X1 U4493 ( .A(n250), .B(n3916), .Y(n3917) );
  CLKINVX1 U4494 ( .A(Input1[74]), .Y(n3916) );
  OAI221X1 U4495 ( .A0(n2200), .A1(n2274), .B0(n3918), .B1(n2273), .C0(n3919), 
        .Y(n1853) );
  MXI2X1 U4496 ( .A(n3920), .B(n3921), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[72]), .Y(n3919) );
  OAI21X1 U4497 ( .A0(n3922), .A1(n282), .B0(n2267), .Y(n3921) );
  NOR2X1 U4498 ( .A(n2082), .B(n2204), .Y(n3922) );
  NOR3X1 U4499 ( .A(n275), .B(n2204), .C(n2082), .Y(n3920) );
  MXI2X1 U4500 ( .A(n3893), .B(n3923), .S0(n308), .Y(n2200) );
  XOR2X1 U4501 ( .A(n3924), .B(n3925), .Y(n3923) );
  XOR2X1 U4502 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .B(n3926), .Y(
        n3925) );
  XOR2X1 U4503 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_19_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .Y(n3893) );
  OAI221X1 U4504 ( .A0(n1490), .A1(n171), .B0(n1854), .B1(n157), .C0(n3927), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_73_N3) );
  AOI22XL U4505 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_73_), 
        .B0(n225), .B1(Input1[73]), .Y(n3927) );
  CLKINVX1 U4506 ( .A(n1491), .Y(n1490) );
  OAI2B2X1 U4507 ( .A1N(Output1[73]), .A0(n2507), .B0(n3928), .B1(n2508), .Y(
        n1491) );
  XNOR2X1 U4508 ( .A(n1854), .B(n3929), .Y(Output1[73]) );
  NOR2X1 U4509 ( .A(n250), .B(n3928), .Y(n3929) );
  CLKINVX1 U4510 ( .A(Input1[73]), .Y(n3928) );
  AOI221XL U4511 ( .A0(n2077), .A1(n2293), .B0(n2082), .B1(n291), .C0(n3930), 
        .Y(n1854) );
  AO22X1 U4512 ( .A0(n267), .A1(n3931), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[75]), .B1(n301), .Y(n3930) );
  CLKINVX1 U4513 ( .A(n3873), .Y(n2077) );
  MXI2X1 U4514 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .B(n3932), .S0(
        n311), .Y(n3873) );
  XOR2X1 U4515 ( .A(n3933), .B(n3934), .Y(n3932) );
  XOR2X1 U4516 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .B(n3935), .Y(
        n3934) );
  OAI221X1 U4517 ( .A0(n1494), .A1(n171), .B0(n1856), .B1(n158), .C0(n3936), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_72_N3) );
  AOI22XL U4518 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_72_), 
        .B0(n225), .B1(Input1[72]), .Y(n3936) );
  CLKINVX1 U4519 ( .A(n1495), .Y(n1494) );
  OAI2B2X1 U4520 ( .A1N(Input1[72]), .A0(n2508), .B0(n3937), .B1(n2507), .Y(
        n1495) );
  CLKNAND2X2 U4521 ( .A(n3836), .B(dec), .Y(n2507) );
  CLKINVX1 U4522 ( .A(Output1[72]), .Y(n3937) );
  XOR2X1 U4523 ( .A(n3938), .B(n1856), .Y(Output1[72]) );
  AOI221XL U4524 ( .A0(n3855), .A1(n297), .B0(n2202), .B1(n2293), .C0(n3939), 
        .Y(n1856) );
  AO22X1 U4525 ( .A0(n267), .A1(n3940), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[72]), .B1(n292), .Y(n3939) );
  CLKINVX1 U4526 ( .A(n3889), .Y(n2202) );
  MXI2X1 U4527 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .B(n3941), .S0(
        n309), .Y(n3889) );
  XOR2X1 U4528 ( .A(n3942), .B(n3943), .Y(n3941) );
  XOR2X1 U4529 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[33]), .B(n3944), .Y(
        n3943) );
  XOR2X1 U4530 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_18_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[72]), .Y(n3855) );
  CLKNAND2X2 U4531 ( .A(Input1[72]), .B(n2288), .Y(n3938) );
  CLKNAND2X2 U4532 ( .A(n3836), .B(n3734), .Y(n2508) );
  OAI221X1 U4533 ( .A0(n3945), .A1(n2300), .B0(n3946), .B1(n2302), .C0(n3947), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_71_N3) );
  AOI22XL U4534 ( .A0(n186), .A1(n1498), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1858), .Y(n3947) );
  OAI222X1 U4535 ( .A0(n2600), .A1(n3948), .B0(n3949), .B1(n3740), .C0(n3946), 
        .C1(n2601), .Y(n1498) );
  CLKINVX1 U4536 ( .A(Output1[71]), .Y(n3948) );
  XOR2X1 U4537 ( .A(n1858), .B(n3950), .Y(Output1[71]) );
  NOR2X1 U4538 ( .A(n250), .B(n3946), .Y(n3950) );
  OAI221X1 U4539 ( .A0(n3951), .A1(n2273), .B0(n2267), .B1(n3952), .C0(n3953), 
        .Y(n1858) );
  AOI222XL U4540 ( .A0(n291), .A1(n2212), .B0(n2258), .B1(n3954), .C0(n2312), 
        .C1(n3955), .Y(n3953) );
  XOR2X1 U4541 ( .A(n3956), .B(n3957), .Y(n3954) );
  XOR2X1 U4542 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[56]), .B(n3958), .Y(
        n3957) );
  CLKINVX1 U4543 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .Y(n3952) );
  CLKINVX1 U4544 ( .A(Input1[71]), .Y(n3946) );
  CLKINVX1 U4545 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_71_), .Y(n3945) );
  OAI221X1 U4546 ( .A0(n1501), .A1(n171), .B0(n1859), .B1(n158), .C0(n3959), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_70_N3) );
  AOI22XL U4547 ( .A0(n197), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_70_), 
        .B0(n225), .B1(Input1[70]), .Y(n3959) );
  CLKINVX1 U4548 ( .A(n1502), .Y(n1501) );
  OAI2B2X1 U4549 ( .A1N(Output1[70]), .A0(n2600), .B0(n3960), .B1(n2601), .Y(
        n1502) );
  CLKINVX1 U4550 ( .A(Input1[70]), .Y(n3960) );
  XOR2X1 U4551 ( .A(n3961), .B(n1859), .Y(Output1[70]) );
  CLKINVX1 U4552 ( .A(n3962), .Y(n1859) );
  OAI221X1 U4553 ( .A0(n3963), .A1(n2274), .B0(n3964), .B1(n2273), .C0(n3965), 
        .Y(n3962) );
  AOI22XL U4554 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[66]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .B1(n291), .Y(n3965) );
  XOR2X1 U4555 ( .A(n3966), .B(n3967), .Y(n3963) );
  MXI2X1 U4556 ( .A(n3968), .B(n3969), .S0(n310), .Y(n3967) );
  XOR2X1 U4557 ( .A(n3970), .B(n3971), .Y(n3969) );
  XNOR2X1 U4558 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .B(n3972), .Y(
        n3970) );
  CLKNAND2X2 U4559 ( .A(n2208), .B(n3973), .Y(n3966) );
  CLKNAND2X2 U4560 ( .A(Input1[70]), .B(n2288), .Y(n3961) );
  OAI221X1 U4561 ( .A0(n3974), .A1(n2300), .B0(n3975), .B1(n2302), .C0(n3976), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_7_N3) );
  AOI22XL U4562 ( .A0(n186), .A1(n1747), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1958), .Y(n3976) );
  CLKINVX1 U4563 ( .A(n1746), .Y(n1747) );
  AOI222XL U4564 ( .A0(n2288), .A1(n3977), .B0(Input1[7]), .B1(n2627), .C0(
        n1989), .C1(Output1[7]), .Y(n1746) );
  XOR2X1 U4565 ( .A(n1958), .B(n3978), .Y(Output1[7]) );
  NOR2X1 U4566 ( .A(n251), .B(n3975), .Y(n3978) );
  OAI221X1 U4567 ( .A0(n3979), .A1(n2273), .B0(n2267), .B1(n3980), .C0(n3981), 
        .Y(n1958) );
  AOI222XL U4568 ( .A0(n291), .A1(n2168), .B0(n2258), .B1(n3982), .C0(n2312), 
        .C1(n3983), .Y(n3981) );
  XOR2X1 U4569 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[8]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[104]), .Y(n3982) );
  CLKINVX1 U4570 ( .A(Input1[7]), .Y(n3975) );
  CLKINVX1 U4571 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_7_), .Y(n3974) );
  OAI221X1 U4572 ( .A0(n1505), .A1(n170), .B0(n3984), .B1(n158), .C0(n3985), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_69_N3) );
  AOI22XL U4573 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_69_), 
        .B0(n225), .B1(Input1[69]), .Y(n3985) );
  CLKINVX1 U4574 ( .A(n1861), .Y(n3984) );
  CLKINVX1 U4575 ( .A(n1506), .Y(n1505) );
  OAI2B2X1 U4576 ( .A1N(Output1[69]), .A0(n2600), .B0(n3986), .B1(n2601), .Y(
        n1506) );
  XOR2X1 U4577 ( .A(n1861), .B(n3987), .Y(Output1[69]) );
  NOR2X1 U4578 ( .A(n251), .B(n3986), .Y(n3987) );
  CLKINVX1 U4579 ( .A(Input1[69]), .Y(n3986) );
  OAI222X1 U4580 ( .A0(n2730), .A1(n3988), .B0(n3989), .B1(n2274), .C0(n3990), 
        .C1(n2273), .Y(n1861) );
  XOR2X1 U4581 ( .A(n3991), .B(n3992), .Y(n3989) );
  MXI2X1 U4582 ( .A(n3993), .B(n3994), .S0(n312), .Y(n3992) );
  XOR2X1 U4583 ( .A(n3995), .B(n3996), .Y(n3994) );
  XNOR2X1 U4584 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .B(n3997), .Y(
        n3995) );
  CLKNAND2X2 U4585 ( .A(n3998), .B(n3999), .Y(n3991) );
  CLKINVX1 U4586 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .Y(n3988) );
  OAI221X1 U4587 ( .A0(n1509), .A1(n170), .B0(n1863), .B1(n157), .C0(n4000), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_68_N3) );
  AOI22XL U4588 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_68_), 
        .B0(n225), .B1(Input1[68]), .Y(n4000) );
  CLKINVX1 U4589 ( .A(n1510), .Y(n1509) );
  OAI2B2X1 U4590 ( .A1N(Input1[68]), .A0(n2601), .B0(n4001), .B1(n2600), .Y(
        n1510) );
  CLKINVX1 U4591 ( .A(Output1[68]), .Y(n4001) );
  XOR2X1 U4592 ( .A(n4002), .B(n1863), .Y(Output1[68]) );
  AOI221XL U4593 ( .A0(n4003), .A1(n297), .B0(n2087), .B1(n2293), .C0(n4004), 
        .Y(n1863) );
  AO22X1 U4594 ( .A0(n266), .A1(n4005), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .B1(n292), .Y(n4004) );
  CLKINVX1 U4595 ( .A(n3998), .Y(n2087) );
  MXI2X1 U4596 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[67]), .B(n4006), .S0(
        n312), .Y(n3998) );
  XOR2X1 U4597 ( .A(n4007), .B(n4008), .Y(n4006) );
  XOR2X1 U4598 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[59]), .B(n4009), .Y(
        n4008) );
  CLKNAND2X2 U4599 ( .A(Input1[68]), .B(n2288), .Y(n4002) );
  OAI221X1 U4600 ( .A0(n1513), .A1(n170), .B0(n4010), .B1(n157), .C0(n4011), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_67_N3) );
  AOI22XL U4601 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_67_), 
        .B0(n225), .B1(Input1[67]), .Y(n4011) );
  CLKINVX1 U4602 ( .A(n1865), .Y(n4010) );
  CLKINVX1 U4603 ( .A(n1514), .Y(n1513) );
  OAI2B2X1 U4604 ( .A1N(Output1[67]), .A0(n2600), .B0(n4012), .B1(n2601), .Y(
        n1514) );
  XOR2X1 U4605 ( .A(n1865), .B(n4013), .Y(Output1[67]) );
  NOR2X1 U4606 ( .A(n251), .B(n4012), .Y(n4013) );
  CLKINVX1 U4607 ( .A(Input1[67]), .Y(n4012) );
  OAI211XL U4608 ( .A0(n4014), .A1(n2273), .B0(n4015), .C0(n4016), .Y(n1865)
         );
  AOI22XL U4609 ( .A0(n2258), .A1(n4017), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[66]), .B1(n2312), .Y(n4016) );
  XNOR2X1 U4610 ( .A(n4018), .B(n4019), .Y(n4017) );
  XOR2X1 U4611 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[58]), .B(n4020), .Y(
        n4019) );
  MXI2X1 U4612 ( .A(n4021), .B(n4022), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[68]), .Y(n4015) );
  OAI21X1 U4613 ( .A0(n4023), .A1(n282), .B0(n2267), .Y(n4022) );
  NOR2X1 U4614 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .Y(n4023) );
  NOR3X1 U4615 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .Y(n4021) );
  OAI221X1 U4616 ( .A0(n1517), .A1(n170), .B0(n4024), .B1(n157), .C0(n4025), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_66_N3) );
  AOI22XL U4617 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_66_), 
        .B0(n225), .B1(Input1[66]), .Y(n4025) );
  CLKINVX1 U4618 ( .A(n1867), .Y(n4024) );
  CLKINVX1 U4619 ( .A(n1518), .Y(n1517) );
  OAI2B2X1 U4620 ( .A1N(Output1[66]), .A0(n2600), .B0(n4026), .B1(n2601), .Y(
        n1518) );
  XOR2X1 U4621 ( .A(n1867), .B(n4027), .Y(Output1[66]) );
  NOR2X1 U4622 ( .A(n251), .B(n4026), .Y(n4027) );
  CLKINVX1 U4623 ( .A(Input1[66]), .Y(n4026) );
  OAI221X1 U4624 ( .A0(n2208), .A1(n2274), .B0(n4028), .B1(n2273), .C0(n4029), 
        .Y(n1867) );
  MXI2X1 U4625 ( .A(n4030), .B(n4031), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[64]), .Y(n4029) );
  OAI21X1 U4626 ( .A0(n4032), .A1(n282), .B0(n2267), .Y(n4031) );
  NOR2X1 U4627 ( .A(n2089), .B(n2212), .Y(n4032) );
  NOR3X1 U4628 ( .A(n275), .B(n2212), .C(n2089), .Y(n4030) );
  MXI2X1 U4629 ( .A(n4003), .B(n4033), .S0(n312), .Y(n2208) );
  XOR2X1 U4630 ( .A(n4034), .B(n4035), .Y(n4033) );
  XOR2X1 U4631 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .B(n4036), .Y(
        n4035) );
  XOR2X1 U4632 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_17_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .Y(n4003) );
  OAI221X1 U4633 ( .A0(n1521), .A1(n170), .B0(n1868), .B1(n157), .C0(n4037), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_65_N3) );
  AOI22XL U4634 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_65_), 
        .B0(n225), .B1(Input1[65]), .Y(n4037) );
  CLKINVX1 U4635 ( .A(n1522), .Y(n1521) );
  OAI2B2X1 U4636 ( .A1N(Output1[65]), .A0(n2600), .B0(n4038), .B1(n2601), .Y(
        n1522) );
  XNOR2X1 U4637 ( .A(n1868), .B(n4039), .Y(Output1[65]) );
  NOR2X1 U4638 ( .A(n251), .B(n4038), .Y(n4039) );
  CLKINVX1 U4639 ( .A(Input1[65]), .Y(n4038) );
  AOI221XL U4640 ( .A0(n2084), .A1(n2293), .B0(n2089), .B1(n291), .C0(n4040), 
        .Y(n1868) );
  AO22X1 U4641 ( .A0(n267), .A1(n4041), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[67]), .B1(n301), .Y(n4040) );
  CLKINVX1 U4642 ( .A(n3973), .Y(n2084) );
  MXI2X1 U4643 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .B(n4042), .S0(
        n312), .Y(n3973) );
  XOR2X1 U4644 ( .A(n4043), .B(n4044), .Y(n4042) );
  XOR2X1 U4645 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .B(n4045), .Y(
        n4044) );
  OAI221X1 U4646 ( .A0(n1525), .A1(n170), .B0(n1870), .B1(n157), .C0(n4046), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_64_N3) );
  AOI22XL U4647 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_64_), 
        .B0(n225), .B1(Input1[64]), .Y(n4046) );
  CLKINVX1 U4648 ( .A(n1526), .Y(n1525) );
  OAI2B2X1 U4649 ( .A1N(Input1[64]), .A0(n2601), .B0(n4047), .B1(n2600), .Y(
        n1526) );
  CLKNAND2X2 U4650 ( .A(n4048), .B(dec), .Y(n2600) );
  CLKINVX1 U4651 ( .A(Output1[64]), .Y(n4047) );
  XOR2X1 U4652 ( .A(n4049), .B(n1870), .Y(Output1[64]) );
  AOI221XL U4653 ( .A0(n3955), .A1(n297), .B0(n2210), .B1(n2293), .C0(n4050), 
        .Y(n1870) );
  AO22X1 U4654 ( .A0(n267), .A1(n4051), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[64]), .B1(n292), .Y(n4050) );
  CLKINVX1 U4655 ( .A(n3999), .Y(n2210) );
  MXI2X1 U4656 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .B(n4052), .S0(
        n312), .Y(n3999) );
  XOR2X1 U4657 ( .A(n4053), .B(n4054), .Y(n4052) );
  XOR2X1 U4658 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[57]), .B(n4055), .Y(
        n4054) );
  XOR2X1 U4659 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_16_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[64]), .Y(n3955) );
  CLKNAND2X2 U4660 ( .A(Input1[64]), .B(n2288), .Y(n4049) );
  CLKNAND2X2 U4661 ( .A(n4048), .B(n3734), .Y(n2601) );
  OA21X1 U4662 ( .A0(Block_Size[0]), .A1(Block_Size[3]), .B0(n3836), .Y(n4048)
         );
  AOI21X1 U4663 ( .A0(n4056), .A1(n4057), .B0(n4058), .Y(n3836) );
  OAI221X1 U4664 ( .A0(n4059), .A1(n2300), .B0(n4060), .B1(n2302), .C0(n4061), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_63_N3) );
  AOI22XL U4665 ( .A0(n186), .A1(n1529), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1872), .Y(n4061) );
  OAI222X1 U4666 ( .A0(n2703), .A1(n4062), .B0(n3628), .B1(n3740), .C0(n4060), 
        .C1(n2704), .Y(n1529) );
  CLKNAND2X2 U4667 ( .A(Block_Size[2]), .B(n4056), .Y(n3740) );
  CLKINVX1 U4668 ( .A(Output1[63]), .Y(n4062) );
  XOR2X1 U4669 ( .A(n1872), .B(n4063), .Y(Output1[63]) );
  NOR2X1 U4670 ( .A(n251), .B(n4060), .Y(n4063) );
  OAI221X1 U4671 ( .A0(n4064), .A1(n277), .B0(n2267), .B1(n4065), .C0(n4066), 
        .Y(n1872) );
  AOI222XL U4672 ( .A0(n2258), .A1(n3747), .B0(n260), .B1(n4067), .C0(n2312), 
        .C1(n4068), .Y(n4066) );
  XOR2X1 U4673 ( .A(n4045), .B(n4069), .Y(n4067) );
  XOR2X1 U4674 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[64]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[40]), .Y(n4069) );
  XOR2X1 U4675 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[39]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_39_), .Y(n4045) );
  XNOR2X1 U4676 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[72]), .B(n3842), .Y(
        n3747) );
  CLKINVX1 U4677 ( .A(Input1[63]), .Y(n4060) );
  CLKINVX1 U4678 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_63_), .Y(n4059) );
  OAI221X1 U4679 ( .A0(n1532), .A1(n170), .B0(n1873), .B1(n157), .C0(n4070), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_62_N3) );
  AOI22XL U4680 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_62_), 
        .B0(n224), .B1(Input1[62]), .Y(n4070) );
  CLKINVX1 U4681 ( .A(n1533), .Y(n1532) );
  OAI2B2X1 U4682 ( .A1N(Output1[62]), .A0(n2703), .B0(n4071), .B1(n2704), .Y(
        n1533) );
  CLKINVX1 U4683 ( .A(Input1[62]), .Y(n4071) );
  XOR2X1 U4684 ( .A(n4072), .B(n1873), .Y(Output1[62]) );
  CLKINVX1 U4685 ( .A(n4073), .Y(n1873) );
  OAI211XL U4686 ( .A0(n285), .A1(n4065), .B0(n4074), .C0(n4075), .Y(n4073) );
  AOI22XL U4687 ( .A0(n262), .A1(n4076), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[58]), .B1(n299), .Y(n4075) );
  XOR2X1 U4688 ( .A(n4036), .B(n4077), .Y(n4076) );
  XOR2X1 U4689 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[68]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .Y(n4077) );
  XOR2X1 U4690 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[38]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_38_), .Y(n4036) );
  MXI2X1 U4691 ( .A(n4078), .B(n4079), .S0(n4080), .Y(n4074) );
  NOR2X1 U4692 ( .A(n2214), .B(n2091), .Y(n4080) );
  CLKINVX1 U4693 ( .A(n4081), .Y(n2091) );
  CLKINVX1 U4694 ( .A(n4082), .Y(n2214) );
  OAI22X1 U4695 ( .A0(n2722), .A1(n3762), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .B1(n2255), .Y(n4079) );
  AO22X1 U4696 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .A1(n2312), .B0(
        n3762), .B1(n2258), .Y(n4078) );
  XNOR2X1 U4697 ( .A(n4083), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[76]), .Y(
        n3762) );
  CLKINVX1 U4698 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[57]), .Y(n4065) );
  CLKNAND2X2 U4699 ( .A(Input1[62]), .B(n2288), .Y(n4072) );
  OAI221X1 U4700 ( .A0(n1536), .A1(n170), .B0(n1874), .B1(n157), .C0(n4084), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_61_N3) );
  AOI22XL U4701 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_61_), 
        .B0(n224), .B1(Input1[61]), .Y(n4084) );
  CLKINVX1 U4702 ( .A(n1537), .Y(n1536) );
  OAI2B2X1 U4703 ( .A1N(Output1[61]), .A0(n2703), .B0(n4085), .B1(n2704), .Y(
        n1537) );
  CLKINVX1 U4704 ( .A(Input1[61]), .Y(n4085) );
  XOR2X1 U4705 ( .A(n4086), .B(n1874), .Y(Output1[61]) );
  CLKINVX1 U4706 ( .A(n4087), .Y(n1874) );
  OAI221X1 U4707 ( .A0(n4088), .A1(n2273), .B0(n2730), .B1(n4089), .C0(n4090), 
        .Y(n4087) );
  MXI2X1 U4708 ( .A(n4091), .B(n4092), .S0(n4093), .Y(n4090) );
  NOR2X1 U4709 ( .A(n2094), .B(n2217), .Y(n4093) );
  OAI22X1 U4710 ( .A0(n2722), .A1(n3777), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .B1(n2255), .Y(n4092) );
  AO22X1 U4711 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .A1(n2312), .B0(
        n3777), .B1(n2258), .Y(n4091) );
  XNOR2X1 U4712 ( .A(n3883), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[8]), .Y(
        n3777) );
  XOR2X1 U4713 ( .A(n4094), .B(n3958), .Y(n4088) );
  XOR2X1 U4714 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[37]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_37_), .Y(n3958) );
  XOR2X1 U4715 ( .A(n3993), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .Y(
        n4094) );
  CLKNAND2X2 U4716 ( .A(Input1[61]), .B(n2288), .Y(n4086) );
  OAI221X1 U4717 ( .A0(n1540), .A1(n170), .B0(n1875), .B1(n157), .C0(n4095), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_60_N3) );
  AOI22XL U4718 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_60_), 
        .B0(n224), .B1(Input1[60]), .Y(n4095) );
  CLKINVX1 U4719 ( .A(n1541), .Y(n1540) );
  OAI2B2X1 U4720 ( .A1N(Output1[60]), .A0(n2703), .B0(n4096), .B1(n2704), .Y(
        n1541) );
  XNOR2X1 U4721 ( .A(n1875), .B(n4097), .Y(Output1[60]) );
  NOR2X1 U4722 ( .A(n251), .B(n4096), .Y(n4097) );
  CLKINVX1 U4723 ( .A(Input1[60]), .Y(n4096) );
  AOI221XL U4724 ( .A0(n2094), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .C0(n4098), .Y(n1875) );
  AO22X1 U4725 ( .A0(n267), .A1(n4099), .B0(n300), .B1(n4100), .Y(n4098) );
  XOR2X1 U4726 ( .A(n2110), .B(n4101), .Y(n4099) );
  XOR2X1 U4727 ( .A(n3972), .B(n2089), .Y(n4101) );
  XOR2X1 U4728 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_17_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[67]), .Y(n2089) );
  XOR2X1 U4729 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[36]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_36_), .Y(n3972) );
  MX2X1 U4730 ( .A(n3788), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[59]), .S0(
        n322), .Y(n2094) );
  XOR2X1 U4731 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[11]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[75]), .Y(n3788) );
  OAI221X1 U4732 ( .A0(n1750), .A1(n170), .B0(n1959), .B1(n157), .C0(n4102), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_6_N3) );
  AOI22XL U4733 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_6_), 
        .B0(n224), .B1(Input1[6]), .Y(n4102) );
  AOI22XL U4734 ( .A0(Input1[6]), .A1(n2627), .B0(n1989), .B1(Output1[6]), .Y(
        n1750) );
  XOR2X1 U4735 ( .A(n4103), .B(n1959), .Y(Output1[6]) );
  CLKINVX1 U4736 ( .A(n4104), .Y(n1959) );
  OAI221X1 U4737 ( .A0(n4105), .A1(n2274), .B0(n4106), .B1(n2273), .C0(n4107), 
        .Y(n4104) );
  AOI22XL U4738 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[2]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[1]), .B1(n291), .Y(n4107) );
  XOR2X1 U4739 ( .A(n4108), .B(n4109), .Y(n4105) );
  MXI2X1 U4740 ( .A(n4110), .B(n4111), .S0(n312), .Y(n4109) );
  XOR2X1 U4741 ( .A(n4112), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[12]), .Y(
        n4111) );
  CLKNAND2X2 U4742 ( .A(n2144), .B(n2025), .Y(n4108) );
  CLKNAND2X2 U4743 ( .A(Input1[6]), .B(n2288), .Y(n4103) );
  OAI221X1 U4744 ( .A0(n1544), .A1(n170), .B0(n4113), .B1(n157), .C0(n4114), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_59_N3) );
  AOI22XL U4745 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_59_), 
        .B0(n224), .B1(Input1[59]), .Y(n4114) );
  CLKINVX1 U4746 ( .A(n1877), .Y(n4113) );
  CLKINVX1 U4747 ( .A(n1545), .Y(n1544) );
  OAI2B2X1 U4748 ( .A1N(Output1[59]), .A0(n2703), .B0(n4115), .B1(n2704), .Y(
        n1545) );
  XOR2X1 U4749 ( .A(n1877), .B(n4116), .Y(Output1[59]) );
  NOR2X1 U4750 ( .A(n251), .B(n4115), .Y(n4116) );
  CLKINVX1 U4751 ( .A(Input1[59]), .Y(n4115) );
  OAI211XL U4752 ( .A0(n3799), .A1(n2722), .B0(n4117), .C0(n4118), .Y(n1877)
         );
  AOI22XL U4753 ( .A0(n262), .A1(n4119), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[58]), .B1(n2312), .Y(n4118) );
  XOR2X1 U4754 ( .A(n4009), .B(n4120), .Y(n4119) );
  XOR2X1 U4755 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[41]), .Y(n4120) );
  XOR2X1 U4756 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[35]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_35_), .Y(n4009) );
  MXI2X1 U4757 ( .A(n4121), .B(n4122), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .Y(n4117) );
  OAI21X1 U4758 ( .A0(n4123), .A1(n282), .B0(n2267), .Y(n4122) );
  NOR2X1 U4759 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .Y(n4123) );
  NOR3X1 U4760 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .Y(n4121) );
  XNOR2X1 U4761 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[74]), .Y(n3799) );
  OAI221X1 U4762 ( .A0(n1548), .A1(n170), .B0(n4124), .B1(n157), .C0(n4125), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_58_N3) );
  AOI22XL U4763 ( .A0(n196), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_58_), 
        .B0(n224), .B1(Input1[58]), .Y(n4125) );
  CLKINVX1 U4764 ( .A(n1879), .Y(n4124) );
  CLKINVX1 U4765 ( .A(n1549), .Y(n1548) );
  OAI2B2X1 U4766 ( .A1N(Output1[58]), .A0(n2703), .B0(n4126), .B1(n2704), .Y(
        n1549) );
  XOR2X1 U4767 ( .A(n1879), .B(n4127), .Y(Output1[58]) );
  NOR2X1 U4768 ( .A(n251), .B(n4126), .Y(n4127) );
  CLKINVX1 U4769 ( .A(Input1[58]), .Y(n4126) );
  OAI221X1 U4770 ( .A0(n4128), .A1(n2273), .B0(n4082), .B1(n2274), .C0(n4129), 
        .Y(n1879) );
  MXI2X1 U4771 ( .A(n4130), .B(n4131), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .Y(n4129) );
  OAI21X1 U4772 ( .A0(n4132), .A1(n282), .B0(n2267), .Y(n4131) );
  NOR2X1 U4773 ( .A(n2219), .B(n2096), .Y(n4132) );
  NOR3X1 U4774 ( .A(n275), .B(n2219), .C(n2096), .Y(n4130) );
  MXI2X1 U4775 ( .A(n4100), .B(n3815), .S0(n312), .Y(n4082) );
  XOR2X1 U4776 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .Y(n3815) );
  XOR2X1 U4777 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_15_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .Y(n4100) );
  XNOR2X1 U4778 ( .A(n4020), .B(n4133), .Y(n4128) );
  XOR2X1 U4779 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .Y(n4133) );
  XOR2X1 U4780 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[34]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_34_), .Y(n4020) );
  OAI221X1 U4781 ( .A0(n1552), .A1(n169), .B0(n1880), .B1(n157), .C0(n4134), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_57_N3) );
  AOI22XL U4782 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_57_), 
        .B0(n224), .B1(Input1[57]), .Y(n4134) );
  CLKINVX1 U4783 ( .A(n1553), .Y(n1552) );
  OAI2B2X1 U4784 ( .A1N(Output1[57]), .A0(n2703), .B0(n4135), .B1(n2704), .Y(
        n1553) );
  CLKINVX1 U4785 ( .A(Input1[57]), .Y(n4135) );
  XOR2X1 U4786 ( .A(n4136), .B(n1880), .Y(Output1[57]) );
  CLKINVX1 U4787 ( .A(n4137), .Y(n1880) );
  OAI221X1 U4788 ( .A0(n4138), .A1(n2273), .B0(n4081), .B1(n2274), .C0(n4139), 
        .Y(n4137) );
  AOI22XL U4789 ( .A0(n291), .A1(n2096), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[59]), .B1(n299), .Y(n4139) );
  MXI2X1 U4790 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .B(n3824), .S0(
        n312), .Y(n4081) );
  XOR2X1 U4791 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .Y(n3824) );
  XNOR2X1 U4792 ( .A(n4055), .B(n4140), .Y(n4138) );
  XOR2X1 U4793 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .Y(n4140) );
  XOR2X1 U4794 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[33]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_33_), .Y(n4055) );
  CLKNAND2X2 U4795 ( .A(Input1[57]), .B(n2288), .Y(n4136) );
  OAI221X1 U4796 ( .A0(n1556), .A1(n169), .B0(n1881), .B1(n157), .C0(n4141), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_56_N3) );
  AOI22XL U4797 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_56_), 
        .B0(n224), .B1(Input1[56]), .Y(n4141) );
  CLKINVX1 U4798 ( .A(n1557), .Y(n1556) );
  OAI2B2X1 U4799 ( .A1N(Output1[56]), .A0(n2703), .B0(n4142), .B1(n2704), .Y(
        n1557) );
  CLKNAND2X2 U4800 ( .A(Block_Size[3]), .B(n3734), .Y(n2704) );
  CLKNAND2X2 U4801 ( .A(dec), .B(Block_Size[3]), .Y(n2703) );
  XNOR2X1 U4802 ( .A(n1881), .B(n4143), .Y(Output1[56]) );
  NOR2X1 U4803 ( .A(n251), .B(n4142), .Y(n4143) );
  CLKINVX1 U4804 ( .A(Input1[56]), .Y(n4142) );
  AOI221XL U4805 ( .A0(n2217), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[56]), .C0(n4144), .Y(n1881) );
  AO22X1 U4806 ( .A0(n267), .A1(n4145), .B0(n301), .B1(n4068), .Y(n4144) );
  XNOR2X1 U4807 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_14_), .B(n4146), .Y(
        n4068) );
  CLKINVX1 U4808 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[56]), .Y(n4146) );
  XOR2X1 U4809 ( .A(n2233), .B(n4147), .Y(n4145) );
  XOR2X1 U4810 ( .A(n2212), .B(n3997), .Y(n4147) );
  XOR2X1 U4811 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[32]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_32_), .Y(n3997) );
  XOR2X1 U4812 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_16_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[66]), .Y(n2212) );
  MX2X1 U4813 ( .A(n3833), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[57]), .S0(
        n322), .Y(n2217) );
  XOR2X1 U4814 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .B(n4148), .Y(
        n3833) );
  OAI221X1 U4815 ( .A0(n4149), .A1(n2300), .B0(n4150), .B1(n2302), .C0(n4151), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_55_N3) );
  AOI22XL U4816 ( .A0(n186), .A1(n1560), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1883), .Y(n4151) );
  OAI222X1 U4817 ( .A0(n2801), .A1(n4152), .B0(n4153), .B1(n4154), .C0(n4150), 
        .C1(n2802), .Y(n1560) );
  CLKINVX1 U4818 ( .A(Output1[55]), .Y(n4152) );
  XOR2X1 U4819 ( .A(n1883), .B(n4155), .Y(Output1[55]) );
  NOR2X1 U4820 ( .A(n251), .B(n4150), .Y(n4155) );
  OAI221X1 U4821 ( .A0(n2267), .A1(n3732), .B0(n4156), .B1(n278), .C0(n4157), 
        .Y(n1883) );
  AOI222XL U4822 ( .A0(n2258), .A1(n3856), .B0(n260), .B1(n4158), .C0(n2312), 
        .C1(n4159), .Y(n4157) );
  XOR2X1 U4823 ( .A(n3722), .B(n4160), .Y(n4158) );
  XOR2X1 U4824 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[88]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[32]), .Y(n4160) );
  XOR2X1 U4825 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[47]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_47_), .Y(n3722) );
  XOR2X1 U4826 ( .A(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[64]), .Y(n3856) );
  CLKINVX1 U4827 ( .A(Input1[55]), .Y(n4150) );
  CLKINVX1 U4828 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_55_), .Y(n4149) );
  OAI221X1 U4829 ( .A0(n1563), .A1(n169), .B0(n1884), .B1(n157), .C0(n4161), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_54_N3) );
  AOI22XL U4830 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_54_), 
        .B0(n224), .B1(Input1[54]), .Y(n4161) );
  CLKINVX1 U4831 ( .A(n1564), .Y(n1563) );
  OAI2B2X1 U4832 ( .A1N(Output1[54]), .A0(n2801), .B0(n4162), .B1(n2802), .Y(
        n1564) );
  CLKINVX1 U4833 ( .A(Input1[54]), .Y(n4162) );
  XOR2X1 U4834 ( .A(n4163), .B(n1884), .Y(Output1[54]) );
  CLKINVX1 U4835 ( .A(n4164), .Y(n1884) );
  AOI22XL U4836 ( .A0(n262), .A1(n4167), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[50]), .B1(n299), .Y(n4166) );
  XOR2X1 U4837 ( .A(n3707), .B(n4168), .Y(n4167) );
  XOR2X1 U4838 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[92]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .Y(n4168) );
  XOR2X1 U4839 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[46]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_46_), .Y(n3707) );
  MXI2X1 U4840 ( .A(n4169), .B(n4170), .S0(n4171), .Y(n4165) );
  NOR2X1 U4841 ( .A(n2221), .B(n2098), .Y(n4171) );
  CLKINVX1 U4842 ( .A(n4172), .Y(n2098) );
  CLKINVX1 U4843 ( .A(n4173), .Y(n2221) );
  OAI22X1 U4844 ( .A0(n2722), .A1(n3871), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[52]), .B1(n2255), .Y(n4170) );
  OAI2BB2X1 U4845 ( .B0(n2255), .B1(n3651), .A0N(n3871), .A1N(n2258), .Y(n4169) );
  XNOR2X1 U4846 ( .A(n4110), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[68]), .Y(
        n3871) );
  CLKINVX1 U4847 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[4]), .Y(n4110) );
  CLKINVX1 U4848 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[52]), .Y(n3651) );
  CLKINVX1 U4849 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[49]), .Y(n3732) );
  CLKNAND2X2 U4850 ( .A(Input1[54]), .B(n2288), .Y(n4163) );
  OAI221X1 U4851 ( .A0(n1567), .A1(n169), .B0(n1885), .B1(n157), .C0(n4174), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_53_N3) );
  AOI22XL U4852 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_53_), 
        .B0(n224), .B1(Input1[53]), .Y(n4174) );
  CLKINVX1 U4853 ( .A(n1568), .Y(n1567) );
  OAI2B2X1 U4854 ( .A1N(Output1[53]), .A0(n2801), .B0(n4175), .B1(n2802), .Y(
        n1568) );
  CLKINVX1 U4855 ( .A(Input1[53]), .Y(n4175) );
  XOR2X1 U4856 ( .A(n4176), .B(n1885), .Y(Output1[53]) );
  CLKINVX1 U4857 ( .A(n4177), .Y(n1885) );
  OAI221X1 U4858 ( .A0(n4178), .A1(n2273), .B0(n2730), .B1(n4179), .C0(n4180), 
        .Y(n4177) );
  MXI2X1 U4859 ( .A(n4181), .B(n4182), .S0(n4183), .Y(n4180) );
  NOR2X1 U4860 ( .A(n2101), .B(n2224), .Y(n4183) );
  OAI22X1 U4861 ( .A0(n2722), .A1(n3886), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .B1(n2255), .Y(n4182) );
  OAI2BB2X1 U4862 ( .B0(n2255), .B1(n4184), .A0N(n3886), .A1N(n2258), .Y(n4181) );
  XNOR2X1 U4863 ( .A(n4185), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[64]), .Y(
        n3886) );
  CLKINVX1 U4864 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .Y(n4184) );
  XOR2X1 U4865 ( .A(n4186), .B(n3637), .Y(n4178) );
  XOR2X1 U4866 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[45]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_45_), .Y(n3637) );
  XOR2X1 U4867 ( .A(n3663), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .Y(
        n4186) );
  CLKINVX1 U4868 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[88]), .Y(n3663) );
  CLKNAND2X2 U4869 ( .A(Input1[53]), .B(n2288), .Y(n4176) );
  OAI221X1 U4870 ( .A0(n1571), .A1(n169), .B0(n1886), .B1(n156), .C0(n4187), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_52_N3) );
  AOI22XL U4871 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_52_), 
        .B0(n224), .B1(Input1[52]), .Y(n4187) );
  CLKINVX1 U4872 ( .A(n1572), .Y(n1571) );
  OAI2B2X1 U4873 ( .A1N(Output1[52]), .A0(n2801), .B0(n4188), .B1(n2802), .Y(
        n1572) );
  XNOR2X1 U4874 ( .A(n1886), .B(n4189), .Y(Output1[52]) );
  NOR2X1 U4875 ( .A(n251), .B(n4188), .Y(n4189) );
  CLKINVX1 U4876 ( .A(Input1[52]), .Y(n4188) );
  AOI221XL U4877 ( .A0(n2101), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .C0(n4190), .Y(n1886) );
  AO22X1 U4878 ( .A0(n267), .A1(n4191), .B0(n301), .B1(n4192), .Y(n4190) );
  XOR2X1 U4879 ( .A(n2117), .B(n4193), .Y(n4191) );
  XOR2X1 U4880 ( .A(n3652), .B(n2068), .Y(n4193) );
  XOR2X1 U4881 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_23_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[91]), .Y(n2068) );
  XOR2X1 U4882 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[44]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_44_), .Y(n3652) );
  MX2X1 U4883 ( .A(n3897), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[51]), .S0(
        n322), .Y(n2101) );
  XOR2X1 U4884 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[3]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[67]), .Y(n3897) );
  OAI221X1 U4885 ( .A0(n1575), .A1(n169), .B0(n4194), .B1(n156), .C0(n4195), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_51_N3) );
  AOI22XL U4886 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_51_), 
        .B0(n224), .B1(Input1[51]), .Y(n4195) );
  CLKINVX1 U4887 ( .A(n1888), .Y(n4194) );
  CLKINVX1 U4888 ( .A(n1576), .Y(n1575) );
  OAI2B2X1 U4889 ( .A1N(Output1[51]), .A0(n2801), .B0(n4196), .B1(n2802), .Y(
        n1576) );
  XOR2X1 U4890 ( .A(n1888), .B(n4197), .Y(Output1[51]) );
  NOR2X1 U4891 ( .A(n251), .B(n4196), .Y(n4197) );
  CLKINVX1 U4892 ( .A(Input1[51]), .Y(n4196) );
  OAI211XL U4893 ( .A0(n3908), .A1(n2722), .B0(n4198), .C0(n4199), .Y(n1888)
         );
  AOI22XL U4894 ( .A0(n262), .A1(n4200), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[50]), .B1(n2312), .Y(n4199) );
  XOR2X1 U4895 ( .A(n3680), .B(n4201), .Y(n4200) );
  XOR2X1 U4896 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[33]), .Y(n4201) );
  XOR2X1 U4897 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[43]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_43_), .Y(n3680) );
  MXI2X1 U4898 ( .A(n4202), .B(n4203), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[52]), .Y(n4198) );
  OAI21X1 U4899 ( .A0(n4204), .A1(n283), .B0(n2267), .Y(n4203) );
  NOR2X1 U4900 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .Y(n4204) );
  NOR3X1 U4901 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .Y(n4202) );
  XNOR2X1 U4902 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[2]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[66]), .Y(n3908) );
  OAI221X1 U4903 ( .A0(n1579), .A1(n169), .B0(n4205), .B1(n156), .C0(n4206), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_50_N3) );
  AOI22XL U4904 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_50_), 
        .B0(n224), .B1(Input1[50]), .Y(n4206) );
  CLKINVX1 U4905 ( .A(n1890), .Y(n4205) );
  CLKINVX1 U4906 ( .A(n1580), .Y(n1579) );
  OAI2B2X1 U4907 ( .A1N(Output1[50]), .A0(n2801), .B0(n4207), .B1(n2802), .Y(
        n1580) );
  XOR2X1 U4908 ( .A(n1890), .B(n4208), .Y(Output1[50]) );
  NOR2X1 U4909 ( .A(n251), .B(n4207), .Y(n4208) );
  CLKINVX1 U4910 ( .A(Input1[50]), .Y(n4207) );
  OAI221X1 U4911 ( .A0(n4209), .A1(n2273), .B0(n4173), .B1(n2274), .C0(n4210), 
        .Y(n1890) );
  MXI2X1 U4912 ( .A(n4211), .B(n4212), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .Y(n4210) );
  OAI21X1 U4913 ( .A0(n4213), .A1(n280), .B0(n2267), .Y(n4212) );
  NOR2X1 U4914 ( .A(n2226), .B(n2103), .Y(n4213) );
  NOR3X1 U4915 ( .A(n276), .B(n2226), .C(n2103), .Y(n4211) );
  MXI2X1 U4916 ( .A(n4192), .B(n3924), .S0(n312), .Y(n4173) );
  XOR2X1 U4917 ( .A(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .Y(n3924) );
  XOR2X1 U4918 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_13_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .Y(n4192) );
  XNOR2X1 U4919 ( .A(n3691), .B(n4214), .Y(n4209) );
  XOR2X1 U4920 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .Y(n4214) );
  XOR2X1 U4921 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[42]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_42_), .Y(n3691) );
  OAI221X1 U4922 ( .A0(n1753), .A1(n169), .B0(n4215), .B1(n156), .C0(n4216), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_5_N3) );
  AOI22XL U4923 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_5_), 
        .B0(n223), .B1(Input1[5]), .Y(n4216) );
  CLKINVX1 U4924 ( .A(n1961), .Y(n4215) );
  AOI22XL U4925 ( .A0(n1989), .A1(Output1[5]), .B0(Input1[5]), .B1(n2627), .Y(
        n1753) );
  XOR2X1 U4926 ( .A(n1961), .B(n4217), .Y(Output1[5]) );
  NOR2BX1 U4927 ( .AN(Input1[5]), .B(n254), .Y(n4217) );
  OAI222X1 U4928 ( .A0(n2730), .A1(n4218), .B0(n4219), .B1(n2274), .C0(n4220), 
        .C1(n2273), .Y(n1961) );
  XOR2X1 U4929 ( .A(n4221), .B(n4222), .Y(n4219) );
  MXI2X1 U4930 ( .A(n4185), .B(n4223), .S0(n312), .Y(n4222) );
  XOR2X1 U4931 ( .A(n4224), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[8]), .Y(
        n4223) );
  CLKNAND2X2 U4932 ( .A(n4225), .B(n4226), .Y(n4221) );
  OAI221X1 U4933 ( .A0(n1583), .A1(n169), .B0(n1891), .B1(n156), .C0(n4227), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_49_N3) );
  AOI22XL U4934 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_49_), 
        .B0(n223), .B1(Input1[49]), .Y(n4227) );
  CLKINVX1 U4935 ( .A(n1584), .Y(n1583) );
  OAI2B2X1 U4936 ( .A1N(Output1[49]), .A0(n2801), .B0(n4228), .B1(n2802), .Y(
        n1584) );
  CLKINVX1 U4937 ( .A(Input1[49]), .Y(n4228) );
  XOR2X1 U4938 ( .A(n4229), .B(n1891), .Y(Output1[49]) );
  CLKINVX1 U4939 ( .A(n4230), .Y(n1891) );
  OAI221X1 U4940 ( .A0(n4231), .A1(n2273), .B0(n4172), .B1(n2274), .C0(n4232), 
        .Y(n4230) );
  AOI22XL U4941 ( .A0(n291), .A1(n2103), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[51]), .B1(n299), .Y(n4232) );
  MXI2X1 U4942 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .B(n3933), .S0(
        n312), .Y(n4172) );
  XOR2X1 U4943 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .Y(n3933) );
  XOR2X1 U4944 ( .A(n4233), .B(n4234), .Y(n4231) );
  XOR2X1 U4945 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .Y(n4234) );
  XOR2X1 U4946 ( .A(n1992), .B(n3733), .Y(n4233) );
  XOR2X1 U4947 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[41]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_41_), .Y(n3733) );
  MXI2X1 U4948 ( .A(n6), .B(n4235), .S0(n1989), .Y(n1992) );
  XOR2X1 U4949 ( .A(Inst_forkAE_CipherInst_CL_n22), .B(
        Inst_forkAE_CipherInst_CL_STATE_0_), .Y(n4235) );
  CLKNAND2X2 U4950 ( .A(Input1[49]), .B(n2288), .Y(n4229) );
  OAI221X1 U4951 ( .A0(n1587), .A1(n169), .B0(n1892), .B1(n156), .C0(n4236), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_48_N3) );
  AOI22XL U4952 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_48_), 
        .B0(n223), .B1(Input1[48]), .Y(n4236) );
  CLKINVX1 U4953 ( .A(n1588), .Y(n1587) );
  OAI2B2X1 U4954 ( .A1N(Output1[48]), .A0(n2801), .B0(n4237), .B1(n2802), .Y(
        n1588) );
  CLKNAND2X2 U4955 ( .A(n4153), .B(n3734), .Y(n2802) );
  CLKNAND2X2 U4956 ( .A(n4153), .B(dec), .Y(n2801) );
  AOI31X1 U4957 ( .A0(n4238), .A1(n4239), .A2(n4057), .B0(n4056), .Y(n4153) );
  XNOR2X1 U4958 ( .A(n1892), .B(n4240), .Y(Output1[48]) );
  NOR2X1 U4959 ( .A(n251), .B(n4237), .Y(n4240) );
  CLKINVX1 U4960 ( .A(Input1[48]), .Y(n4237) );
  AOI221XL U4961 ( .A0(n2224), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[48]), .C0(n4241), .Y(n1892) );
  AO22X1 U4962 ( .A0(n267), .A1(n4242), .B0(n301), .B1(n4159), .Y(n4241) );
  XNOR2X1 U4963 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_12_), .B(n4243), .Y(
        n4159) );
  CLKINVX1 U4964 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[48]), .Y(n4243) );
  XOR2X1 U4965 ( .A(n4244), .B(n4245), .Y(n4242) );
  XOR2X1 U4966 ( .A(n1991), .B(n2240), .Y(n4245) );
  MXI2X1 U4967 ( .A(n461), .B(n4), .S0(n1989), .Y(n1991) );
  XNOR2X1 U4968 ( .A(n3667), .B(n2188), .Y(n4244) );
  XOR2X1 U4969 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_22_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[90]), .Y(n2188) );
  XOR2X1 U4970 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[40]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_40_), .Y(n3667) );
  MX2X1 U4971 ( .A(n3942), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[49]), .S0(
        n321), .Y(n2224) );
  XOR2X1 U4972 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[1]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .Y(n3942) );
  OAI221X1 U4973 ( .A0(n4246), .A1(n2300), .B0(n4247), .B1(n2302), .C0(n4248), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_47_N3) );
  AOI22XL U4974 ( .A0(n186), .A1(n1591), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1894), .Y(n4248) );
  OAI222X1 U4975 ( .A0(n2894), .A1(n4249), .B0(n3849), .B1(n4154), .C0(n4247), 
        .C1(n2895), .Y(n1591) );
  CLKINVX1 U4976 ( .A(Output1[47]), .Y(n4249) );
  XOR2X1 U4977 ( .A(n1894), .B(n4250), .Y(Output1[47]) );
  NOR2X1 U4978 ( .A(n252), .B(n4247), .Y(n4250) );
  OAI221X1 U4979 ( .A0(n4251), .A1(n277), .B0(n2267), .B1(n4252), .C0(n4253), 
        .Y(n1894) );
  AOI222XL U4980 ( .A0(n2258), .A1(n3956), .B0(n260), .B1(n4254), .C0(n2312), 
        .C1(n4255), .Y(n4253) );
  XOR2X1 U4981 ( .A(n3826), .B(n4256), .Y(n4254) );
  XOR2X1 U4982 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[80]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[56]), .Y(n4256) );
  XOR2X1 U4983 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[15]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_15_), .Y(n3826) );
  XOR2X1 U4984 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[24]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[88]), .Y(n3956) );
  CLKINVX1 U4985 ( .A(Input1[47]), .Y(n4247) );
  CLKINVX1 U4986 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_47_), .Y(n4246) );
  OAI221X1 U4987 ( .A0(n1594), .A1(n169), .B0(n1895), .B1(n156), .C0(n4257), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_46_N3) );
  AOI22XL U4988 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_46_), 
        .B0(n223), .B1(Input1[46]), .Y(n4257) );
  CLKINVX1 U4989 ( .A(n1595), .Y(n1594) );
  OAI2B2X1 U4990 ( .A1N(Output1[46]), .A0(n2894), .B0(n4258), .B1(n2895), .Y(
        n1595) );
  CLKINVX1 U4991 ( .A(Input1[46]), .Y(n4258) );
  XOR2X1 U4992 ( .A(n4259), .B(n1895), .Y(Output1[46]) );
  CLKINVX1 U4993 ( .A(n4260), .Y(n1895) );
  OAI211XL U4994 ( .A0(n285), .A1(n4252), .B0(n4261), .C0(n4262), .Y(n4260) );
  AOI22XL U4995 ( .A0(n261), .A1(n4263), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[42]), .B1(n299), .Y(n4262) );
  XOR2X1 U4996 ( .A(n3817), .B(n4264), .Y(n4263) );
  XOR2X1 U4997 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[84]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .Y(n4264) );
  XOR2X1 U4998 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[14]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_14_), .Y(n3817) );
  MXI2X1 U4999 ( .A(n4265), .B(n4266), .S0(n4267), .Y(n4261) );
  NOR2X1 U5000 ( .A(n2228), .B(n2105), .Y(n4267) );
  CLKINVX1 U5001 ( .A(n4268), .Y(n2105) );
  CLKINVX1 U5002 ( .A(n4269), .Y(n2228) );
  OAI22X1 U5003 ( .A0(n2722), .A1(n3971), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .B1(n2255), .Y(n4266) );
  AO22X1 U5004 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .A1(n2312), .B0(
        n3971), .B1(n2258), .Y(n4265) );
  XNOR2X1 U5005 ( .A(n4270), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[92]), .Y(
        n3971) );
  CLKINVX1 U5006 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[41]), .Y(n4252) );
  CLKNAND2X2 U5007 ( .A(Input1[46]), .B(n2288), .Y(n4259) );
  OAI221X1 U5008 ( .A0(n1598), .A1(n169), .B0(n1896), .B1(n156), .C0(n4271), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_45_N3) );
  AOI22XL U5009 ( .A0(n195), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_45_), 
        .B0(n223), .B1(Input1[45]), .Y(n4271) );
  CLKINVX1 U5010 ( .A(n1599), .Y(n1598) );
  OAI2B2X1 U5011 ( .A1N(Output1[45]), .A0(n2894), .B0(n4272), .B1(n2895), .Y(
        n1599) );
  CLKINVX1 U5012 ( .A(Input1[45]), .Y(n4272) );
  XOR2X1 U5013 ( .A(n4273), .B(n1896), .Y(Output1[45]) );
  CLKINVX1 U5014 ( .A(n4274), .Y(n1896) );
  OAI221X1 U5015 ( .A0(n4275), .A1(n2273), .B0(n2730), .B1(n4276), .C0(n4277), 
        .Y(n4274) );
  MXI2X1 U5016 ( .A(n4278), .B(n4279), .S0(n4280), .Y(n4277) );
  NOR2X1 U5017 ( .A(n2108), .B(n2231), .Y(n4280) );
  OAI22X1 U5018 ( .A0(n2722), .A1(n3996), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .B1(n2255), .Y(n4279) );
  AO22X1 U5019 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .A1(n2312), .B0(
        n3996), .B1(n2258), .Y(n4278) );
  XNOR2X1 U5020 ( .A(n4281), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[88]), .Y(
        n3996) );
  XOR2X1 U5021 ( .A(n4282), .B(n3749), .Y(n4275) );
  XOR2X1 U5022 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[13]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_13_), .Y(n3749) );
  XOR2X1 U5023 ( .A(n3774), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .Y(
        n4282) );
  CLKNAND2X2 U5024 ( .A(Input1[45]), .B(n2288), .Y(n4273) );
  OAI221X1 U5025 ( .A0(n1602), .A1(n168), .B0(n1897), .B1(n156), .C0(n4283), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_44_N3) );
  AOI22XL U5026 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_44_), 
        .B0(n223), .B1(Input1[44]), .Y(n4283) );
  CLKINVX1 U5027 ( .A(n1603), .Y(n1602) );
  OAI2B2X1 U5028 ( .A1N(Output1[44]), .A0(n2894), .B0(n4284), .B1(n2895), .Y(
        n1603) );
  XNOR2X1 U5029 ( .A(n1897), .B(n4285), .Y(Output1[44]) );
  NOR2X1 U5030 ( .A(n252), .B(n4284), .Y(n4285) );
  CLKINVX1 U5031 ( .A(Input1[44]), .Y(n4284) );
  AOI221XL U5032 ( .A0(n2108), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .C0(n4286), .Y(n1897) );
  AO22X1 U5033 ( .A0(n267), .A1(n4287), .B0(n300), .B1(n4288), .Y(n4286) );
  XOR2X1 U5034 ( .A(n2096), .B(n4289), .Y(n4287) );
  XOR2X1 U5035 ( .A(n3763), .B(n2075), .Y(n4289) );
  XOR2X1 U5036 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_21_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[83]), .Y(n2075) );
  XOR2X1 U5037 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[12]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_12_), .Y(n3763) );
  MX2X1 U5038 ( .A(n4007), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[43]), .S0(
        n320), .Y(n2108) );
  XOR2X1 U5039 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[27]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[91]), .Y(n4007) );
  OAI221X1 U5040 ( .A0(n1606), .A1(n168), .B0(n4290), .B1(n156), .C0(n4291), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_43_N3) );
  AOI22XL U5041 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_43_), 
        .B0(n223), .B1(Input1[43]), .Y(n4291) );
  CLKINVX1 U5042 ( .A(n1899), .Y(n4290) );
  CLKINVX1 U5043 ( .A(n1607), .Y(n1606) );
  OAI2B2X1 U5044 ( .A1N(Output1[43]), .A0(n2894), .B0(n4292), .B1(n2895), .Y(
        n1607) );
  XOR2X1 U5045 ( .A(n1899), .B(n4293), .Y(Output1[43]) );
  NOR2X1 U5046 ( .A(n252), .B(n4292), .Y(n4293) );
  CLKINVX1 U5047 ( .A(Input1[43]), .Y(n4292) );
  OAI211XL U5048 ( .A0(n4018), .A1(n2722), .B0(n4294), .C0(n4295), .Y(n1899)
         );
  AOI22XL U5049 ( .A0(n262), .A1(n4296), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[42]), .B1(n2312), .Y(n4295) );
  XOR2X1 U5050 ( .A(n3790), .B(n4297), .Y(n4296) );
  XOR2X1 U5051 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[57]), .Y(n4297) );
  XOR2X1 U5052 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[11]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_11_), .Y(n3790) );
  MXI2X1 U5053 ( .A(n4298), .B(n4299), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .Y(n4294) );
  OAI21X1 U5054 ( .A0(n4300), .A1(n281), .B0(n2267), .Y(n4299) );
  NOR2X1 U5055 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .Y(n4300) );
  NOR3X1 U5056 ( .A(n285), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .Y(n4298) );
  XNOR2X1 U5057 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[26]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[90]), .Y(n4018) );
  OAI221X1 U5058 ( .A0(n1610), .A1(n168), .B0(n4301), .B1(n156), .C0(n4302), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_42_N3) );
  AOI22XL U5059 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_42_), 
        .B0(n223), .B1(Input1[42]), .Y(n4302) );
  CLKINVX1 U5060 ( .A(n1901), .Y(n4301) );
  CLKINVX1 U5061 ( .A(n1611), .Y(n1610) );
  OAI2B2X1 U5062 ( .A1N(Output1[42]), .A0(n2894), .B0(n4303), .B1(n2895), .Y(
        n1611) );
  XOR2X1 U5063 ( .A(n1901), .B(n4304), .Y(Output1[42]) );
  NOR2X1 U5064 ( .A(n252), .B(n4303), .Y(n4304) );
  CLKINVX1 U5065 ( .A(Input1[42]), .Y(n4303) );
  OAI221X1 U5066 ( .A0(n4305), .A1(n2273), .B0(n4269), .B1(n2274), .C0(n4306), 
        .Y(n1901) );
  MXI2X1 U5067 ( .A(n4307), .B(n4308), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .Y(n4306) );
  OAI21X1 U5068 ( .A0(n4309), .A1(n283), .B0(n2267), .Y(n4308) );
  NOR2X1 U5069 ( .A(n2110), .B(n2233), .Y(n4309) );
  NOR3X1 U5070 ( .A(n278), .B(n2110), .C(n2233), .Y(n4307) );
  CLKINVX1 U5071 ( .A(n4251), .Y(n2233) );
  MXI2X1 U5072 ( .A(n4288), .B(n4034), .S0(n312), .Y(n4269) );
  XOR2X1 U5073 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .Y(n4034) );
  XOR2X1 U5074 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_11_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .Y(n4288) );
  XNOR2X1 U5075 ( .A(n3801), .B(n4310), .Y(n4305) );
  XOR2X1 U5076 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .Y(n4310) );
  XNOR2X1 U5077 ( .A(n4311), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_10_), 
        .Y(n3801) );
  OAI221X1 U5078 ( .A0(n1614), .A1(n168), .B0(n1902), .B1(n156), .C0(n4312), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_41_N3) );
  AOI22XL U5079 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_41_), 
        .B0(n223), .B1(Input1[41]), .Y(n4312) );
  CLKINVX1 U5080 ( .A(n1615), .Y(n1614) );
  OAI2B2X1 U5081 ( .A1N(Output1[41]), .A0(n2894), .B0(n4313), .B1(n2895), .Y(
        n1615) );
  CLKINVX1 U5082 ( .A(Input1[41]), .Y(n4313) );
  XOR2X1 U5083 ( .A(n4314), .B(n1902), .Y(Output1[41]) );
  CLKINVX1 U5084 ( .A(n4315), .Y(n1902) );
  OAI221X1 U5085 ( .A0(n2273), .A1(n4316), .B0(n4268), .B1(n2274), .C0(n4317), 
        .Y(n4315) );
  AOI22XL U5086 ( .A0(n291), .A1(n2110), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[43]), .B1(n299), .Y(n4317) );
  MXI2X1 U5087 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .B(n4043), .S0(
        n313), .Y(n4268) );
  XOR2X1 U5088 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .Y(n4043) );
  XOR2X1 U5089 ( .A(n3835), .B(n4318), .Y(n4316) );
  XOR2X1 U5090 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .Y(n4318) );
  XOR2X1 U5091 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[9]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_9_), .Y(n3835) );
  CLKNAND2X2 U5092 ( .A(Input1[41]), .B(n2288), .Y(n4314) );
  OAI221X1 U5093 ( .A0(n1618), .A1(n168), .B0(n1903), .B1(n156), .C0(n4319), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_40_N3) );
  AOI22XL U5094 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_40_), 
        .B0(n223), .B1(Input1[40]), .Y(n4319) );
  CLKINVX1 U5095 ( .A(n1619), .Y(n1618) );
  OAI2B2X1 U5096 ( .A1N(Output1[40]), .A0(n2894), .B0(n4320), .B1(n2895), .Y(
        n1619) );
  CLKNAND2X2 U5097 ( .A(n4321), .B(n3734), .Y(n2895) );
  CLKNAND2X2 U5098 ( .A(dec), .B(n4321), .Y(n2894) );
  OAI21X1 U5099 ( .A0(n4056), .A1(n4057), .B0(n4322), .Y(n4321) );
  XNOR2X1 U5100 ( .A(n1903), .B(n4323), .Y(Output1[40]) );
  NOR2X1 U5101 ( .A(n252), .B(n4320), .Y(n4323) );
  CLKINVX1 U5102 ( .A(Input1[40]), .Y(n4320) );
  AOI221XL U5103 ( .A0(n2231), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[40]), .C0(n4324), .Y(n1903) );
  AO22X1 U5104 ( .A0(n267), .A1(n4325), .B0(n300), .B1(n4255), .Y(n4324) );
  XNOR2X1 U5105 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_10_), .B(n4326), .Y(
        n4255) );
  CLKINVX1 U5106 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[40]), .Y(n4326) );
  XOR2X1 U5107 ( .A(n3778), .B(n4327), .Y(n4325) );
  XOR2X1 U5108 ( .A(n2219), .B(n2196), .Y(n4327) );
  XOR2X1 U5109 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_20_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[82]), .Y(n2196) );
  XOR2X1 U5110 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[8]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_8_), .Y(n3778) );
  MX2X1 U5111 ( .A(n4053), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[41]), .S0(
        n319), .Y(n2231) );
  XOR2X1 U5112 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[25]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .Y(n4053) );
  OAI221X1 U5113 ( .A0(n1756), .A1(n168), .B0(n1963), .B1(n156), .C0(n4328), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_4_N3) );
  AOI22XL U5114 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_4_), 
        .B0(n223), .B1(Input1[4]), .Y(n4328) );
  AOI22XL U5115 ( .A0(Input1[4]), .A1(n2627), .B0(n1989), .B1(Output1[4]), .Y(
        n1756) );
  XOR2X1 U5116 ( .A(n4329), .B(n1963), .Y(Output1[4]) );
  AOI221XL U5117 ( .A0(n4330), .A1(n297), .B0(n2047), .B1(n2293), .C0(n4331), 
        .Y(n1963) );
  AO22X1 U5118 ( .A0(n268), .A1(n4332), .B0(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .B1(n292), .Y(n4331) );
  CLKINVX1 U5119 ( .A(n4225), .Y(n2047) );
  MXI2X1 U5120 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[3]), .B(n4333), .S0(
        n313), .Y(n4225) );
  XOR2X1 U5121 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[11]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[107]), .Y(n4333) );
  CLKNAND2X2 U5122 ( .A(Input1[4]), .B(n2288), .Y(n4329) );
  OAI221X1 U5123 ( .A0(n4334), .A1(n2300), .B0(n4335), .B1(n2302), .C0(n4336), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_39_N3) );
  AOI22XL U5124 ( .A0(n186), .A1(n1622), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1905), .Y(n4336) );
  OAI222X1 U5125 ( .A0(n2984), .A1(n4337), .B0(n3949), .B1(n4154), .C0(n4335), 
        .C1(n2985), .Y(n1622) );
  CLKINVX1 U5126 ( .A(Output1[39]), .Y(n4337) );
  XOR2X1 U5127 ( .A(n1905), .B(n4338), .Y(Output1[39]) );
  NOR2X1 U5128 ( .A(n252), .B(n4335), .Y(n4338) );
  OAI221X1 U5129 ( .A0(n4339), .A1(n277), .B0(n2267), .B1(n4340), .C0(n4341), 
        .Y(n1905) );
  AOI222XL U5130 ( .A0(n2258), .A1(n3635), .B0(n260), .B1(n4342), .C0(n2312), 
        .C1(n4343), .Y(n4341) );
  XOR2X1 U5131 ( .A(n3935), .B(n4344), .Y(n4342) );
  XOR2X1 U5132 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[72]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[48]), .Y(n4344) );
  XOR2X1 U5133 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[31]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_31_), .Y(n3935) );
  XOR2X1 U5134 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[16]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[80]), .Y(n3635) );
  CLKINVX1 U5135 ( .A(Input1[39]), .Y(n4335) );
  CLKINVX1 U5136 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_39_), .Y(n4334) );
  OAI221X1 U5137 ( .A0(n1625), .A1(n168), .B0(n1906), .B1(n156), .C0(n4345), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_38_N3) );
  AOI22XL U5138 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_38_), 
        .B0(n223), .B1(Input1[38]), .Y(n4345) );
  CLKINVX1 U5139 ( .A(n1626), .Y(n1625) );
  OAI2B2X1 U5140 ( .A1N(Output1[38]), .A0(n2984), .B0(n4346), .B1(n2985), .Y(
        n1626) );
  CLKINVX1 U5141 ( .A(Input1[38]), .Y(n4346) );
  XOR2X1 U5142 ( .A(n4347), .B(n1906), .Y(Output1[38]) );
  CLKINVX1 U5143 ( .A(n4348), .Y(n1906) );
  OAI211XL U5144 ( .A0(n285), .A1(n4340), .B0(n4349), .C0(n4350), .Y(n4348) );
  AOI22XL U5145 ( .A0(n262), .A1(n4351), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[34]), .B1(n299), .Y(n4350) );
  XOR2X1 U5146 ( .A(n3926), .B(n4352), .Y(n4351) );
  XOR2X1 U5147 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[76]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[52]), .Y(n4352) );
  XOR2X1 U5148 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[30]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_30_), .Y(n3926) );
  MXI2X1 U5149 ( .A(n4353), .B(n4354), .S0(n4355), .Y(n4349) );
  NOR2X1 U5150 ( .A(n2235), .B(n2112), .Y(n4355) );
  CLKINVX1 U5151 ( .A(n4356), .Y(n2112) );
  CLKINVX1 U5152 ( .A(n4357), .Y(n2235) );
  OAI22X1 U5153 ( .A0(n2722), .A1(n3650), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .B1(n2255), .Y(n4354) );
  AO22X1 U5154 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .A1(n2312), .B0(
        n3650), .B1(n2258), .Y(n4353) );
  XNOR2X1 U5155 ( .A(n4358), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[84]), .Y(
        n3650) );
  CLKINVX1 U5156 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[33]), .Y(n4340) );
  CLKNAND2X2 U5157 ( .A(Input1[38]), .B(n2288), .Y(n4347) );
  OAI221X1 U5158 ( .A0(n1629), .A1(n168), .B0(n1907), .B1(n155), .C0(n4359), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_37_N3) );
  AOI22XL U5159 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_37_), 
        .B0(n223), .B1(Input1[37]), .Y(n4359) );
  CLKINVX1 U5160 ( .A(n1630), .Y(n1629) );
  OAI2B2X1 U5161 ( .A1N(Output1[37]), .A0(n2984), .B0(n4360), .B1(n2985), .Y(
        n1630) );
  CLKINVX1 U5162 ( .A(Input1[37]), .Y(n4360) );
  XOR2X1 U5163 ( .A(n4361), .B(n1907), .Y(Output1[37]) );
  CLKINVX1 U5164 ( .A(n4362), .Y(n1907) );
  OAI221X1 U5165 ( .A0(n4363), .A1(n2273), .B0(n2730), .B1(n4364), .C0(n4365), 
        .Y(n4362) );
  MXI2X1 U5166 ( .A(n4366), .B(n4367), .S0(n4368), .Y(n4365) );
  NOR2X1 U5167 ( .A(n2115), .B(n2238), .Y(n4368) );
  OAI22X1 U5168 ( .A0(n2722), .A1(n3668), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .B1(n2255), .Y(n4367) );
  AO22X1 U5169 ( .A0(n3668), .A1(n2258), .B0(n2312), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .Y(n4366) );
  XOR2X1 U5170 ( .A(n4369), .B(n3774), .Y(n3668) );
  CLKINVX1 U5171 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .Y(n4364) );
  XOR2X1 U5172 ( .A(n4370), .B(n3858), .Y(n4363) );
  XOR2X1 U5173 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[29]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_29_), .Y(n3858) );
  XOR2X1 U5174 ( .A(n3883), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .Y(
        n4370) );
  CLKNAND2X2 U5175 ( .A(Input1[37]), .B(n2288), .Y(n4361) );
  OAI221X1 U5176 ( .A0(n1633), .A1(n168), .B0(n1908), .B1(n155), .C0(n4371), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_36_N3) );
  AOI22XL U5177 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_36_), 
        .B0(n222), .B1(Input1[36]), .Y(n4371) );
  CLKINVX1 U5178 ( .A(n1634), .Y(n1633) );
  OAI2B2X1 U5179 ( .A1N(Output1[36]), .A0(n2984), .B0(n4372), .B1(n2985), .Y(
        n1634) );
  XNOR2X1 U5180 ( .A(n1908), .B(n4373), .Y(Output1[36]) );
  NOR2X1 U5181 ( .A(n252), .B(n4372), .Y(n4373) );
  CLKINVX1 U5182 ( .A(Input1[36]), .Y(n4372) );
  AOI221XL U5183 ( .A0(n2115), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .C0(n4374), .Y(n1908) );
  AO22X1 U5184 ( .A0(n268), .A1(n4375), .B0(n300), .B1(n4376), .Y(n4374) );
  XOR2X1 U5185 ( .A(n2103), .B(n4377), .Y(n4375) );
  XOR2X1 U5186 ( .A(n3872), .B(n2082), .Y(n4377) );
  XOR2X1 U5187 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_19_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[75]), .Y(n2082) );
  XOR2X1 U5188 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[28]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_28_), .Y(n3872) );
  MX2X1 U5189 ( .A(n3678), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[35]), .S0(
        n318), .Y(n2115) );
  XOR2X1 U5190 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[19]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[83]), .Y(n3678) );
  OAI221X1 U5191 ( .A0(n1637), .A1(n168), .B0(n4378), .B1(n155), .C0(n4379), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_35_N3) );
  AOI22XL U5192 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_35_), 
        .B0(n222), .B1(Input1[35]), .Y(n4379) );
  CLKINVX1 U5193 ( .A(n1910), .Y(n4378) );
  CLKINVX1 U5194 ( .A(n1638), .Y(n1637) );
  OAI2B2X1 U5195 ( .A1N(Output1[35]), .A0(n2984), .B0(n4380), .B1(n2985), .Y(
        n1638) );
  XOR2X1 U5196 ( .A(n1910), .B(n4381), .Y(Output1[35]) );
  NOR2X1 U5197 ( .A(n252), .B(n4380), .Y(n4381) );
  CLKINVX1 U5198 ( .A(Input1[35]), .Y(n4380) );
  OAI211XL U5199 ( .A0(n3689), .A1(n2722), .B0(n4382), .C0(n4383), .Y(n1910)
         );
  AOI22XL U5200 ( .A0(n261), .A1(n4384), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[34]), .B1(n2312), .Y(n4383) );
  XOR2X1 U5201 ( .A(n3899), .B(n4385), .Y(n4384) );
  XOR2X1 U5202 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[49]), .Y(n4385) );
  XOR2X1 U5203 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[27]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_27_), .Y(n3899) );
  MXI2X1 U5204 ( .A(n4386), .B(n4387), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .Y(n4382) );
  OAI21X1 U5205 ( .A0(n4388), .A1(n283), .B0(n2267), .Y(n4387) );
  NOR2X1 U5206 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .Y(n4388) );
  NOR3X1 U5207 ( .A(n2266), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .Y(n4386) );
  XNOR2X1 U5208 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[18]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[82]), .Y(n3689) );
  OAI221X1 U5209 ( .A0(n1641), .A1(n168), .B0(n4389), .B1(n155), .C0(n4390), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_34_N3) );
  AOI22XL U5210 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_34_), 
        .B0(n222), .B1(Input1[34]), .Y(n4390) );
  CLKINVX1 U5211 ( .A(n1912), .Y(n4389) );
  CLKINVX1 U5212 ( .A(n1642), .Y(n1641) );
  OAI2B2X1 U5213 ( .A1N(Output1[34]), .A0(n2984), .B0(n4391), .B1(n2985), .Y(
        n1642) );
  XOR2X1 U5214 ( .A(n1912), .B(n4392), .Y(Output1[34]) );
  NOR2X1 U5215 ( .A(n252), .B(n4391), .Y(n4392) );
  CLKINVX1 U5216 ( .A(Input1[34]), .Y(n4391) );
  OAI221X1 U5217 ( .A0(n4393), .A1(n2273), .B0(n4357), .B1(n2274), .C0(n4394), 
        .Y(n1912) );
  MXI2X1 U5218 ( .A(n4395), .B(n4396), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .Y(n4394) );
  OAI21X1 U5219 ( .A0(n4397), .A1(n282), .B0(n2267), .Y(n4396) );
  NOR2X1 U5220 ( .A(n2117), .B(n2240), .Y(n4397) );
  NOR3X1 U5221 ( .A(n279), .B(n2117), .C(n2240), .Y(n4395) );
  CLKINVX1 U5222 ( .A(n4339), .Y(n2240) );
  MXI2X1 U5223 ( .A(n4376), .B(n3705), .S0(n313), .Y(n4357) );
  XOR2X1 U5224 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .Y(n3705) );
  XOR2X1 U5225 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_9_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .Y(n4376) );
  XNOR2X1 U5226 ( .A(n3910), .B(n4398), .Y(n4393) );
  XOR2X1 U5227 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .Y(n4398) );
  XOR2X1 U5228 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[26]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_26_), .Y(n3910) );
  OAI221X1 U5229 ( .A0(n1645), .A1(n168), .B0(n1913), .B1(n155), .C0(n4399), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_33_N3) );
  AOI22XL U5230 ( .A0(n194), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_33_), 
        .B0(n222), .B1(Input1[33]), .Y(n4399) );
  CLKINVX1 U5231 ( .A(n1646), .Y(n1645) );
  OAI2B2X1 U5232 ( .A1N(Output1[33]), .A0(n2984), .B0(n4400), .B1(n2985), .Y(
        n1646) );
  CLKINVX1 U5233 ( .A(Input1[33]), .Y(n4400) );
  XOR2X1 U5234 ( .A(n4401), .B(n1913), .Y(Output1[33]) );
  CLKINVX1 U5235 ( .A(n4402), .Y(n1913) );
  OAI221X1 U5236 ( .A0(n4403), .A1(n2273), .B0(n4356), .B1(n2274), .C0(n4404), 
        .Y(n4402) );
  AOI22XL U5237 ( .A0(n291), .A1(n2117), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[35]), .B1(n299), .Y(n4404) );
  MXI2X1 U5238 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .B(n3720), .S0(
        n313), .Y(n4356) );
  XOR2X1 U5239 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .Y(n3720) );
  XNOR2X1 U5240 ( .A(n3944), .B(n4405), .Y(n4403) );
  XOR2X1 U5241 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .Y(n4405) );
  XOR2X1 U5242 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[25]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_25_), .Y(n3944) );
  CLKNAND2X2 U5243 ( .A(Input1[33]), .B(n2288), .Y(n4401) );
  OAI221X1 U5244 ( .A0(n1649), .A1(n167), .B0(n1914), .B1(n155), .C0(n4406), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_32_N3) );
  AOI22XL U5245 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_32_), 
        .B0(n222), .B1(Input1[32]), .Y(n4406) );
  CLKINVX1 U5246 ( .A(n1650), .Y(n1649) );
  OAI2B2X1 U5247 ( .A1N(Output1[32]), .A0(n2984), .B0(n4407), .B1(n2985), .Y(
        n1650) );
  CLKNAND2X2 U5248 ( .A(n4408), .B(n3734), .Y(n2985) );
  CLKNAND2X2 U5249 ( .A(dec), .B(n4408), .Y(n2984) );
  OAI21X1 U5250 ( .A0(n4056), .A1(n3628), .B0(n4322), .Y(n4408) );
  XNOR2X1 U5251 ( .A(n1914), .B(n4409), .Y(Output1[32]) );
  NOR2X1 U5252 ( .A(n252), .B(n4407), .Y(n4409) );
  CLKINVX1 U5253 ( .A(Input1[32]), .Y(n4407) );
  AOI221XL U5254 ( .A0(n2238), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[32]), .C0(n4410), .Y(n1914) );
  AO22X1 U5255 ( .A0(n268), .A1(n4411), .B0(n300), .B1(n4343), .Y(n4410) );
  XNOR2X1 U5256 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_8_), .B(n4412), .Y(
        n4343) );
  CLKINVX1 U5257 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[32]), .Y(n4412) );
  XOR2X1 U5258 ( .A(n3887), .B(n4413), .Y(n4411) );
  XOR2X1 U5259 ( .A(n2226), .B(n2204), .Y(n4413) );
  XOR2X1 U5260 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_18_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[74]), .Y(n2204) );
  XOR2X1 U5261 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[24]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_24_), .Y(n3887) );
  MX2X1 U5262 ( .A(n3731), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[33]), .S0(
        n317), .Y(n2238) );
  XOR2X1 U5263 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[17]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .Y(n3731) );
  OAI221X1 U5264 ( .A0(n4414), .A1(n2300), .B0(n4415), .B1(n2302), .C0(n4416), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_31_N3) );
  AOI22XL U5265 ( .A0(n186), .A1(n1653), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1916), .Y(n4416) );
  OAI222X1 U5266 ( .A0(n3068), .A1(n4417), .B0(n3628), .B1(n4154), .C0(n4415), 
        .C1(n3069), .Y(n1653) );
  CLKNAND2X2 U5267 ( .A(Block_Size[3]), .B(n4239), .Y(n4154) );
  CLKNAND2X2 U5268 ( .A(Block_Size[0]), .B(Block_Size[1]), .Y(n3628) );
  CLKINVX1 U5269 ( .A(Output1[31]), .Y(n4417) );
  XOR2X1 U5270 ( .A(n1916), .B(n4418), .Y(Output1[31]) );
  NOR2X1 U5271 ( .A(n252), .B(n4415), .Y(n4418) );
  OAI221X1 U5272 ( .A0(n4419), .A1(n2273), .B0(n2267), .B1(n3591), .C0(n4420), 
        .Y(n1916) );
  AOI222XL U5273 ( .A0(n291), .A1(n2124), .B0(n2258), .B1(n4421), .C0(n2312), 
        .C1(n4422), .Y(n4420) );
  XOR2X1 U5274 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[96]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]), .Y(n4421) );
  CLKINVX1 U5275 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[25]), .Y(n3591) );
  CLKINVX1 U5276 ( .A(Input1[31]), .Y(n4415) );
  CLKINVX1 U5277 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_31_), .Y(n4414) );
  OAI221X1 U5278 ( .A0(n1656), .A1(n167), .B0(n1917), .B1(n155), .C0(n4423), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_30_N3) );
  AOI22XL U5279 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_30_), 
        .B0(n222), .B1(Input1[30]), .Y(n4423) );
  CLKINVX1 U5280 ( .A(n1657), .Y(n1656) );
  OAI2B2X1 U5281 ( .A1N(Output1[30]), .A0(n3068), .B0(n4424), .B1(n3069), .Y(
        n1657) );
  CLKINVX1 U5282 ( .A(Input1[30]), .Y(n4424) );
  XOR2X1 U5283 ( .A(n4425), .B(n1917), .Y(Output1[30]) );
  CLKINVX1 U5284 ( .A(n4426), .Y(n1917) );
  OAI221X1 U5285 ( .A0(n4427), .A1(n2274), .B0(n4428), .B1(n2273), .C0(n4429), 
        .Y(n4426) );
  AOI22XL U5286 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[26]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[25]), .B1(n291), .Y(n4429) );
  XOR2X1 U5287 ( .A(n4430), .B(n4431), .Y(n4427) );
  MXI2X1 U5288 ( .A(n4270), .B(n4432), .S0(n313), .Y(n4431) );
  XOR2X1 U5289 ( .A(n4433), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[4]), .Y(
        n4432) );
  CLKINVX1 U5290 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[28]), .Y(n4270) );
  CLKNAND2X2 U5291 ( .A(n2245), .B(n4434), .Y(n4430) );
  CLKNAND2X2 U5292 ( .A(Input1[30]), .B(n2288), .Y(n4425) );
  OAI221X1 U5293 ( .A0(n1759), .A1(n167), .B0(n4435), .B1(n155), .C0(n4436), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_3_N3) );
  AOI22XL U5294 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_3_), 
        .B0(n222), .B1(Input1[3]), .Y(n4436) );
  CLKINVX1 U5295 ( .A(n1965), .Y(n4435) );
  AOI22XL U5296 ( .A0(n1989), .A1(Output1[3]), .B0(Input1[3]), .B1(n2627), .Y(
        n1759) );
  XOR2X1 U5297 ( .A(n1965), .B(n4437), .Y(Output1[3]) );
  NOR2BX1 U5298 ( .AN(Input1[3]), .B(n254), .Y(n4437) );
  OAI211XL U5299 ( .A0(n3592), .A1(n2273), .B0(n4438), .C0(n4439), .Y(n1965)
         );
  AOI22XL U5300 ( .A0(n2258), .A1(n4440), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[2]), .B1(n2312), .Y(n4439) );
  XOR2X1 U5301 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[106]), .Y(n4440) );
  MXI2X1 U5302 ( .A(n4441), .B(n4442), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[4]), .Y(n4438) );
  OAI21X1 U5303 ( .A0(n4443), .A1(n283), .B0(n2267), .Y(n4442) );
  NOR2X1 U5304 ( .A(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .Y(n4443) );
  NOR3X1 U5305 ( .A(n283), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .C(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .Y(n4441) );
  XOR2X1 U5306 ( .A(n4014), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[49]), .Y(
        n3592) );
  XOR2X1 U5307 ( .A(n4444), .B(n4445), .Y(n4014) );
  OAI221X1 U5308 ( .A0(n1660), .A1(n167), .B0(n4446), .B1(n155), .C0(n4447), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_29_N3) );
  AOI22XL U5309 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_29_), 
        .B0(n222), .B1(Input1[29]), .Y(n4447) );
  CLKINVX1 U5310 ( .A(n1919), .Y(n4446) );
  CLKINVX1 U5311 ( .A(n1661), .Y(n1660) );
  OAI2B2X1 U5312 ( .A1N(Output1[29]), .A0(n3068), .B0(n4448), .B1(n3069), .Y(
        n1661) );
  XOR2X1 U5313 ( .A(n1919), .B(n4449), .Y(Output1[29]) );
  NOR2X1 U5314 ( .A(n252), .B(n4448), .Y(n4449) );
  CLKINVX1 U5315 ( .A(Input1[29]), .Y(n4448) );
  OAI222X1 U5316 ( .A0(n2730), .A1(n4450), .B0(n4451), .B1(n2274), .C0(n4452), 
        .C1(n2273), .Y(n1919) );
  XOR2X1 U5317 ( .A(n4453), .B(n4454), .Y(n4451) );
  MXI2X1 U5318 ( .A(n4281), .B(n4455), .S0(n313), .Y(n4454) );
  XOR2X1 U5319 ( .A(n4185), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[96]), .Y(
        n4455) );
  CLKNAND2X2 U5320 ( .A(n4456), .B(n4457), .Y(n4453) );
  CLKINVX1 U5321 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .Y(n4450) );
  OAI221X1 U5322 ( .A0(n1664), .A1(n167), .B0(n1921), .B1(n155), .C0(n4458), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_28_N3) );
  AOI22XL U5323 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_28_), 
        .B0(n222), .B1(Input1[28]), .Y(n4458) );
  CLKINVX1 U5324 ( .A(n1665), .Y(n1664) );
  OAI2B2X1 U5325 ( .A1N(Input1[28]), .A0(n3069), .B0(n4459), .B1(n3068), .Y(
        n1665) );
  CLKINVX1 U5326 ( .A(Output1[28]), .Y(n4459) );
  XOR2X1 U5327 ( .A(n4460), .B(n1921), .Y(Output1[28]) );
  AOI221XL U5328 ( .A0(n4461), .A1(n297), .B0(n2004), .B1(n2293), .C0(n4462), 
        .Y(n1921) );
  OAI2BB2X1 U5329 ( .B0(n4463), .B1(n284), .A0N(n4464), .A1N(n269), .Y(n4462)
         );
  CLKINVX1 U5330 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .Y(n4463) );
  CLKINVX1 U5331 ( .A(n4456), .Y(n2004) );
  MXI2X1 U5332 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[27]), .B(n4465), .S0(
        n313), .Y(n4456) );
  XOR2X1 U5333 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[99]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[3]), .Y(n4465) );
  CLKNAND2X2 U5334 ( .A(Input1[28]), .B(n2288), .Y(n4460) );
  OAI221X1 U5335 ( .A0(n1668), .A1(n167), .B0(n4466), .B1(n155), .C0(n4467), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_27_N3) );
  AOI22XL U5336 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_27_), 
        .B0(n222), .B1(Input1[27]), .Y(n4467) );
  CLKINVX1 U5337 ( .A(n1923), .Y(n4466) );
  CLKINVX1 U5338 ( .A(n1669), .Y(n1668) );
  OAI2B2X1 U5339 ( .A1N(Output1[27]), .A0(n3068), .B0(n4468), .B1(n3069), .Y(
        n1669) );
  XOR2X1 U5340 ( .A(n1923), .B(n4469), .Y(Output1[27]) );
  NOR2X1 U5341 ( .A(n252), .B(n4468), .Y(n4469) );
  CLKINVX1 U5342 ( .A(Input1[27]), .Y(n4468) );
  OAI211XL U5343 ( .A0(n4470), .A1(n2273), .B0(n4471), .C0(n4472), .Y(n1923)
         );
  AOI22XL U5344 ( .A0(n2258), .A1(n4473), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[26]), .B1(n2312), .Y(n4472) );
  XOR2X1 U5345 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[98]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[2]), .Y(n4473) );
  MXI2X1 U5346 ( .A(n4474), .B(n4475), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[28]), .Y(n4471) );
  OAI21X1 U5347 ( .A0(n4476), .A1(n283), .B0(n2267), .Y(n4475) );
  NOR2X1 U5348 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .Y(n4476) );
  NOR3X1 U5349 ( .A(n275), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .Y(n4474) );
  OAI221X1 U5350 ( .A0(n1672), .A1(n167), .B0(n4477), .B1(n155), .C0(n4478), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_26_N3) );
  AOI22XL U5351 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_26_), 
        .B0(n222), .B1(Input1[26]), .Y(n4478) );
  CLKINVX1 U5352 ( .A(n1925), .Y(n4477) );
  CLKINVX1 U5353 ( .A(n1673), .Y(n1672) );
  OAI2B2X1 U5354 ( .A1N(Output1[26]), .A0(n3068), .B0(n4479), .B1(n3069), .Y(
        n1673) );
  XOR2X1 U5355 ( .A(n1925), .B(n4480), .Y(Output1[26]) );
  NOR2X1 U5356 ( .A(n253), .B(n4479), .Y(n4480) );
  CLKINVX1 U5357 ( .A(Input1[26]), .Y(n4479) );
  OAI221X1 U5358 ( .A0(n2245), .A1(n2274), .B0(n4481), .B1(n2273), .C0(n4482), 
        .Y(n1925) );
  MXI2X1 U5359 ( .A(n4483), .B(n4484), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[24]), .Y(n4482) );
  OAI21X1 U5360 ( .A0(n4485), .A1(n283), .B0(n2267), .Y(n4484) );
  NOR2X1 U5361 ( .A(n2124), .B(n2007), .Y(n4485) );
  NOR3X1 U5362 ( .A(n281), .B(n2124), .C(n2007), .Y(n4483) );
  XOR2X1 U5363 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_6_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[26]), .Y(n2124) );
  MXI2X1 U5364 ( .A(n4461), .B(n4486), .S0(n313), .Y(n2245) );
  XOR2X1 U5365 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .B(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .Y(n4486) );
  XOR2X1 U5366 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_7_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .Y(n4461) );
  OAI221X1 U5367 ( .A0(n1676), .A1(n167), .B0(n1927), .B1(n155), .C0(n4487), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_25_N3) );
  AOI22XL U5368 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_25_), 
        .B0(n222), .B1(Input1[25]), .Y(n4487) );
  CLKINVX1 U5369 ( .A(n1677), .Y(n1676) );
  OAI2B2X1 U5370 ( .A1N(Input1[25]), .A0(n3069), .B0(n4488), .B1(n3068), .Y(
        n1677) );
  CLKINVX1 U5371 ( .A(Output1[25]), .Y(n4488) );
  XOR2X1 U5372 ( .A(n4489), .B(n1927), .Y(Output1[25]) );
  AOI221XL U5373 ( .A0(n2119), .A1(n2293), .B0(n261), .B1(n4490), .C0(n4491), 
        .Y(n1927) );
  AO22X1 U5374 ( .A0(n292), .A1(n2007), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[27]), .B1(n302), .Y(n4491) );
  CLKINVX1 U5375 ( .A(n4434), .Y(n2119) );
  MXI2X1 U5376 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .B(n4492), .S0(
        n313), .Y(n4434) );
  XOR2X1 U5377 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .Y(n4492) );
  CLKNAND2X2 U5378 ( .A(Input1[25]), .B(n2288), .Y(n4489) );
  OAI221X1 U5379 ( .A0(n1680), .A1(n167), .B0(n1929), .B1(n155), .C0(n4493), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_24_N3) );
  AOI22XL U5380 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_24_), 
        .B0(n222), .B1(Input1[24]), .Y(n4493) );
  CLKINVX1 U5381 ( .A(n1681), .Y(n1680) );
  OAI2B2X1 U5382 ( .A1N(Input1[24]), .A0(n3069), .B0(n4494), .B1(n3068), .Y(
        n1681) );
  CLKNAND2X2 U5383 ( .A(dec), .B(n4495), .Y(n3068) );
  CLKINVX1 U5384 ( .A(Output1[24]), .Y(n4494) );
  XOR2X1 U5385 ( .A(n4496), .B(n1929), .Y(Output1[24]) );
  AOI221XL U5386 ( .A0(n4422), .A1(n297), .B0(n2122), .B1(n2293), .C0(n4497), 
        .Y(n1929) );
  OAI2BB2X1 U5387 ( .B0(n4498), .B1(n284), .A0N(n4499), .A1N(n269), .Y(n4497)
         );
  CLKINVX1 U5388 ( .A(n4457), .Y(n2122) );
  MXI2X1 U5389 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[25]), .B(n4500), .S0(
        n313), .Y(n4457) );
  XOR2X1 U5390 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[97]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[1]), .Y(n4500) );
  XOR2X1 U5391 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_6_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[24]), .Y(n4422) );
  CLKNAND2X2 U5392 ( .A(Input1[24]), .B(n2288), .Y(n4496) );
  CLKNAND2X2 U5393 ( .A(n4495), .B(n3734), .Y(n3069) );
  OAI221X1 U5394 ( .A0(n4501), .A1(n2300), .B0(n4502), .B1(n2302), .C0(n4503), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_23_N3) );
  AOI22XL U5395 ( .A0(n186), .A1(n1684), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1931), .Y(n4503) );
  OAI222X1 U5396 ( .A0(n4502), .A1(n3153), .B0(n3152), .B1(n4504), .C0(n4322), 
        .C1(n4505), .Y(n1684) );
  CLKINVX1 U5397 ( .A(Output1[23]), .Y(n4504) );
  XOR2X1 U5398 ( .A(n1931), .B(n4506), .Y(Output1[23]) );
  NOR2X1 U5399 ( .A(n253), .B(n4502), .Y(n4506) );
  OAI221X1 U5400 ( .A0(n4507), .A1(n2273), .B0(n2267), .B1(n4508), .C0(n4509), 
        .Y(n1931) );
  AOI222XL U5401 ( .A0(n291), .A1(n2132), .B0(n2258), .B1(n4510), .C0(n2312), 
        .C1(n4511), .Y(n4509) );
  XOR2X1 U5402 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[24]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[120]), .Y(n4510) );
  CLKINVX1 U5403 ( .A(Input1[23]), .Y(n4502) );
  CLKINVX1 U5404 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_23_), .Y(n4501) );
  OAI221X1 U5405 ( .A0(n1687), .A1(n167), .B0(n1932), .B1(n155), .C0(n4512), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_22_N3) );
  AOI22XL U5406 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_22_), 
        .B0(n221), .B1(Input1[22]), .Y(n4512) );
  CLKINVX1 U5407 ( .A(n1688), .Y(n1687) );
  OAI2B2X1 U5408 ( .A1N(Output1[22]), .A0(n3152), .B0(n4513), .B1(n3153), .Y(
        n1688) );
  CLKINVX1 U5409 ( .A(Input1[22]), .Y(n4513) );
  XOR2X1 U5410 ( .A(n4514), .B(n1932), .Y(Output1[22]) );
  CLKINVX1 U5411 ( .A(n4515), .Y(n1932) );
  OAI221X1 U5412 ( .A0(n4516), .A1(n2274), .B0(n4517), .B1(n2273), .C0(n4518), 
        .Y(n4515) );
  AOI22XL U5413 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[18]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[17]), .B1(n292), .Y(n4518) );
  XOR2X1 U5414 ( .A(n4519), .B(n4520), .Y(n4516) );
  MXI2X1 U5415 ( .A(n4358), .B(n4521), .S0(n313), .Y(n4520) );
  XOR2X1 U5416 ( .A(n4522), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[28]), .Y(
        n4521) );
  CLKINVX1 U5417 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[20]), .Y(n4358) );
  CLKNAND2X2 U5418 ( .A(n2128), .B(n4523), .Y(n4519) );
  CLKNAND2X2 U5419 ( .A(Input1[22]), .B(n2288), .Y(n4514) );
  OAI221X1 U5420 ( .A0(n1691), .A1(n167), .B0(n1933), .B1(n155), .C0(n4524), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_21_N3) );
  AOI22XL U5421 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_21_), 
        .B0(n221), .B1(Input1[21]), .Y(n4524) );
  CLKINVX1 U5422 ( .A(n1692), .Y(n1691) );
  OAI2B2X1 U5423 ( .A1N(Output1[21]), .A0(n3152), .B0(n4525), .B1(n3153), .Y(
        n1692) );
  XNOR2X1 U5424 ( .A(n1933), .B(n4526), .Y(Output1[21]) );
  NOR2X1 U5425 ( .A(n252), .B(n4525), .Y(n4526) );
  CLKINVX1 U5426 ( .A(Input1[21]), .Y(n4525) );
  AOI222XL U5427 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), 
        .B0(n4527), .B1(n2293), .C0(n4528), .C1(n265), .Y(n1933) );
  XNOR2X1 U5428 ( .A(n4529), .B(n4530), .Y(n4527) );
  MXI2X1 U5429 ( .A(n4369), .B(n4531), .S0(n313), .Y(n4530) );
  XOR2X1 U5430 ( .A(n4532), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[24]), .Y(
        n4531) );
  CLKINVX1 U5431 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[16]), .Y(n4369) );
  CLKNAND2X2 U5432 ( .A(n4533), .B(n4534), .Y(n4529) );
  OAI221X1 U5433 ( .A0(n1695), .A1(n167), .B0(n1935), .B1(n154), .C0(n4535), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_20_N3) );
  AOI22XL U5434 ( .A0(n193), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_20_), 
        .B0(n221), .B1(Input1[20]), .Y(n4535) );
  CLKINVX1 U5435 ( .A(n1696), .Y(n1695) );
  OAI2B2X1 U5436 ( .A1N(Input1[20]), .A0(n3153), .B0(n4536), .B1(n3152), .Y(
        n1696) );
  CLKINVX1 U5437 ( .A(Output1[20]), .Y(n4536) );
  XOR2X1 U5438 ( .A(n4537), .B(n1935), .Y(Output1[20]) );
  AOI221XL U5439 ( .A0(n4538), .A1(n297), .B0(n2012), .B1(n2293), .C0(n4539), 
        .Y(n1935) );
  AO22X1 U5440 ( .A0(n268), .A1(n4540), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .B1(n292), .Y(n4539) );
  CLKINVX1 U5441 ( .A(n4533), .Y(n2012) );
  MXI2X1 U5442 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[19]), .B(n4541), .S0(
        n314), .Y(n4533) );
  XOR2X1 U5443 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[27]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[123]), .Y(n4541) );
  CLKNAND2X2 U5444 ( .A(Input1[20]), .B(n2288), .Y(n4537) );
  OAI221X1 U5445 ( .A0(n1762), .A1(n166), .B0(n4542), .B1(n154), .C0(n4543), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_2_N3) );
  AOI22XL U5446 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_2_), 
        .B0(n221), .B1(Input1[2]), .Y(n4543) );
  CLKINVX1 U5447 ( .A(n1967), .Y(n4542) );
  AOI22XL U5448 ( .A0(n1989), .A1(Output1[2]), .B0(Input1[2]), .B1(n2627), .Y(
        n1762) );
  XOR2X1 U5449 ( .A(n1967), .B(n4544), .Y(Output1[2]) );
  NOR2BX1 U5450 ( .AN(Input1[2]), .B(n254), .Y(n4544) );
  OAI221X1 U5451 ( .A0(n2144), .A1(n2274), .B0(n3607), .B1(n2273), .C0(n4545), 
        .Y(n1967) );
  MXI2X1 U5452 ( .A(n4546), .B(n4547), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[0]), .Y(n4545) );
  OAI21X1 U5453 ( .A0(n4548), .A1(n283), .B0(n2267), .Y(n4547) );
  NOR2X1 U5454 ( .A(n2049), .B(n2168), .Y(n4548) );
  NOR3X1 U5455 ( .A(n2266), .B(n2168), .C(n2049), .Y(n4546) );
  XOR2X1 U5456 ( .A(n4028), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[52]), .Y(
        n3607) );
  XNOR2X1 U5457 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .B(n3593), .Y(
        n4028) );
  XOR2X1 U5458 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[18]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_18_), .Y(n3593) );
  MXI2X1 U5459 ( .A(n4330), .B(n4549), .S0(n314), .Y(n2144) );
  XOR2X1 U5460 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .Y(n4549) );
  XOR2X1 U5461 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_1_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .Y(n4330) );
  OAI221X1 U5462 ( .A0(n1699), .A1(n166), .B0(n4550), .B1(n154), .C0(n4551), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_19_N3) );
  AOI22XL U5463 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_19_), 
        .B0(n221), .B1(Input1[19]), .Y(n4551) );
  CLKINVX1 U5464 ( .A(n1937), .Y(n4550) );
  CLKINVX1 U5465 ( .A(n1700), .Y(n1699) );
  OAI2B2X1 U5466 ( .A1N(Output1[19]), .A0(n3152), .B0(n4552), .B1(n3153), .Y(
        n1700) );
  XOR2X1 U5467 ( .A(n1937), .B(n4553), .Y(Output1[19]) );
  NOR2X1 U5468 ( .A(n253), .B(n4552), .Y(n4553) );
  CLKINVX1 U5469 ( .A(Input1[19]), .Y(n4552) );
  OAI211XL U5470 ( .A0(n4554), .A1(n2273), .B0(n4555), .C0(n4556), .Y(n1937)
         );
  AOI22XL U5471 ( .A0(n2258), .A1(n4557), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[18]), .B1(n2312), .Y(n4556) );
  XOR2X1 U5472 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[26]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[122]), .Y(n4557) );
  MXI2X1 U5473 ( .A(n4558), .B(n4559), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[20]), .Y(n4555) );
  OAI21X1 U5474 ( .A0(n4560), .A1(n282), .B0(n2267), .Y(n4559) );
  NOR2X1 U5475 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .Y(n4560) );
  NOR3X1 U5476 ( .A(n2266), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .Y(n4558) );
  OAI221X1 U5477 ( .A0(n1703), .A1(n166), .B0(n4561), .B1(n154), .C0(n4562), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_18_N3) );
  AOI22XL U5478 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_18_), 
        .B0(n221), .B1(Input1[18]), .Y(n4562) );
  CLKINVX1 U5479 ( .A(n1939), .Y(n4561) );
  CLKINVX1 U5480 ( .A(n1704), .Y(n1703) );
  OAI2B2X1 U5481 ( .A1N(Output1[18]), .A0(n3152), .B0(n4563), .B1(n3153), .Y(
        n1704) );
  XOR2X1 U5482 ( .A(n1939), .B(n4564), .Y(Output1[18]) );
  NOR2X1 U5483 ( .A(n252), .B(n4563), .Y(n4564) );
  CLKINVX1 U5484 ( .A(Input1[18]), .Y(n4563) );
  OAI221X1 U5485 ( .A0(n2128), .A1(n2274), .B0(n4565), .B1(n2273), .C0(n4566), 
        .Y(n1939) );
  MXI2X1 U5486 ( .A(n4567), .B(n4568), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[16]), .Y(n4566) );
  OAI21X1 U5487 ( .A0(n4569), .A1(n283), .B0(n2267), .Y(n4568) );
  NOR2X1 U5488 ( .A(n2014), .B(n2132), .Y(n4569) );
  NOR3X1 U5489 ( .A(n2266), .B(n2132), .C(n2014), .Y(n4567) );
  MXI2X1 U5490 ( .A(n4538), .B(n4570), .S0(n314), .Y(n2128) );
  XOR2X1 U5491 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[28]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .Y(n4570) );
  XOR2X1 U5492 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_5_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .Y(n4538) );
  OAI221X1 U5493 ( .A0(n1707), .A1(n166), .B0(n1940), .B1(n154), .C0(n4571), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_17_N3) );
  AOI22XL U5494 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_17_), 
        .B0(n221), .B1(Input1[17]), .Y(n4571) );
  CLKINVX1 U5495 ( .A(n1708), .Y(n1707) );
  OAI2B2X1 U5496 ( .A1N(Output1[17]), .A0(n3152), .B0(n4572), .B1(n3153), .Y(
        n1708) );
  XNOR2X1 U5497 ( .A(n1940), .B(n4573), .Y(Output1[17]) );
  NOR2X1 U5498 ( .A(n253), .B(n4572), .Y(n4573) );
  CLKINVX1 U5499 ( .A(Input1[17]), .Y(n4572) );
  AOI221XL U5500 ( .A0(n2009), .A1(n2293), .B0(n2014), .B1(n291), .C0(n4574), 
        .Y(n1940) );
  AO22X1 U5501 ( .A0(n268), .A1(n4575), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[19]), .B1(n302), .Y(n4574) );
  CLKINVX1 U5502 ( .A(n4523), .Y(n2009) );
  MXI2X1 U5503 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .B(n4576), .S0(
        n314), .Y(n4523) );
  XOR2X1 U5504 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[31]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .Y(n4576) );
  OAI221X1 U5505 ( .A0(n1711), .A1(n166), .B0(n1942), .B1(n154), .C0(n4577), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_16_N3) );
  AOI22XL U5506 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_16_), 
        .B0(n221), .B1(Input1[16]), .Y(n4577) );
  CLKINVX1 U5507 ( .A(n1712), .Y(n1711) );
  OAI2B2X1 U5508 ( .A1N(Input1[16]), .A0(n3153), .B0(n4578), .B1(n3152), .Y(
        n1712) );
  CLKNAND2X2 U5509 ( .A(dec), .B(n4505), .Y(n3152) );
  CLKINVX1 U5510 ( .A(Output1[16]), .Y(n4578) );
  XOR2X1 U5511 ( .A(n4579), .B(n1942), .Y(Output1[16]) );
  AOI221XL U5512 ( .A0(n4511), .A1(n297), .B0(n2130), .B1(n2293), .C0(n4580), 
        .Y(n1942) );
  OAI2BB2X1 U5513 ( .B0(n4581), .B1(n285), .A0N(n4582), .A1N(n269), .Y(n4580)
         );
  CLKINVX1 U5514 ( .A(n4534), .Y(n2130) );
  MXI2X1 U5515 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[17]), .B(n4583), .S0(
        n314), .Y(n4534) );
  XOR2X1 U5516 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[25]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[121]), .Y(n4583) );
  XOR2X1 U5517 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_4_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[16]), .Y(n4511) );
  CLKNAND2X2 U5518 ( .A(Input1[16]), .B(n2288), .Y(n4579) );
  CLKNAND2X2 U5519 ( .A(n4505), .B(n3734), .Y(n3153) );
  OAI21X1 U5520 ( .A0(n4322), .A1(n4238), .B0(n4584), .Y(n4505) );
  OAI221X1 U5521 ( .A0(n4585), .A1(n2300), .B0(n4586), .B1(n2302), .C0(n4587), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_15_N3) );
  AOI22XL U5522 ( .A0(n186), .A1(n1715), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1944), .Y(n4587) );
  OAI222X1 U5523 ( .A0(n2379), .A1(n4588), .B0(n4322), .B1(n3849), .C0(n4586), 
        .C1(n2381), .Y(n1715) );
  CLKNAND2X2 U5524 ( .A(Block_Size[0]), .B(n4057), .Y(n3849) );
  CLKINVX1 U5525 ( .A(Output1[15]), .Y(n4588) );
  XOR2X1 U5526 ( .A(n1944), .B(n4589), .Y(Output1[15]) );
  NOR2X1 U5527 ( .A(n253), .B(n4586), .Y(n4589) );
  OAI221X1 U5528 ( .A0(n4590), .A1(n277), .B0(n2267), .B1(n4148), .C0(n4591), 
        .Y(n1944) );
  AOI222XL U5529 ( .A0(n260), .A1(n4592), .B0(n2258), .B1(n4593), .C0(n2312), 
        .C1(n3840), .Y(n4591) );
  XOR2X1 U5530 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_2_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[8]), .Y(n3840) );
  XOR2X1 U5531 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[16]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[112]), .Y(n4593) );
  CLKINVX1 U5532 ( .A(Input1[15]), .Y(n4586) );
  CLKINVX1 U5533 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_15_), .Y(n4585) );
  OAI221X1 U5534 ( .A0(n1718), .A1(n166), .B0(n1945), .B1(n154), .C0(n4594), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_14_N3) );
  AOI22XL U5535 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_14_), 
        .B0(n221), .B1(Input1[14]), .Y(n4594) );
  CLKINVX1 U5536 ( .A(n1719), .Y(n1718) );
  OAI2B2X1 U5537 ( .A1N(Output1[14]), .A0(n2379), .B0(n4595), .B1(n2381), .Y(
        n1719) );
  CLKINVX1 U5538 ( .A(Input1[14]), .Y(n4595) );
  XOR2X1 U5539 ( .A(n4596), .B(n1945), .Y(Output1[14]) );
  CLKINVX1 U5540 ( .A(n4597), .Y(n1945) );
  OAI221X1 U5541 ( .A0(n4598), .A1(n2274), .B0(n4599), .B1(n2273), .C0(n4600), 
        .Y(n4597) );
  AOI22XL U5542 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[10]), .A1(n298), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[9]), .B1(n292), .Y(n4600) );
  XOR2X1 U5543 ( .A(n4601), .B(n4602), .Y(n4598) );
  MXI2X1 U5544 ( .A(n4083), .B(n4603), .S0(n314), .Y(n4602) );
  XOR2X1 U5545 ( .A(n4604), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[20]), .Y(
        n4603) );
  CLKINVX1 U5546 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[12]), .Y(n4083) );
  CLKNAND2X2 U5547 ( .A(n3713), .B(n2136), .Y(n4601) );
  MXI2X1 U5548 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .B(n4605), .S0(
        n314), .Y(n3713) );
  XOR2X1 U5549 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .Y(n4605) );
  CLKNAND2X2 U5550 ( .A(Input1[14]), .B(n2288), .Y(n4596) );
  OAI221X1 U5551 ( .A0(n1722), .A1(n166), .B0(n1946), .B1(n154), .C0(n4606), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_13_N3) );
  AOI22XL U5552 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_13_), 
        .B0(n221), .B1(Input1[13]), .Y(n4606) );
  CLKINVX1 U5553 ( .A(n1723), .Y(n1722) );
  OAI2B2X1 U5554 ( .A1N(Output1[13]), .A0(n2379), .B0(n4607), .B1(n2381), .Y(
        n1723) );
  XNOR2X1 U5555 ( .A(n1946), .B(n4608), .Y(Output1[13]) );
  NOR2X1 U5556 ( .A(n253), .B(n4607), .Y(n4608) );
  CLKINVX1 U5557 ( .A(Input1[13]), .Y(n4607) );
  AOI222XL U5558 ( .A0(n2332), .A1(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), 
        .B0(n4609), .B1(n2293), .C0(n4610), .C1(n265), .Y(n1946) );
  XNOR2X1 U5559 ( .A(n4611), .B(n4612), .Y(n4609) );
  MXI2X1 U5560 ( .A(n4613), .B(n4614), .S0(n314), .Y(n4612) );
  XOR2X1 U5561 ( .A(n4615), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[16]), .Y(
        n4614) );
  CLKNAND2X2 U5562 ( .A(n3844), .B(n4616), .Y(n4611) );
  MXI2X1 U5563 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[9]), .B(n4617), .S0(
        n314), .Y(n3844) );
  XOR2X1 U5564 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[17]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[113]), .Y(n4617) );
  OAI221X1 U5565 ( .A0(n4618), .A1(n2300), .B0(n4619), .B1(n2302), .C0(n4620), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_127_N3) );
  AOI2BB2X1 U5566 ( .B0(n182), .B1(n1288), .A0N(n159), .A1N(n1772), .Y(n4620)
         );
  CLKINVX1 U5567 ( .A(n1287), .Y(n1288) );
  MXI2X1 U5568 ( .A(Input1[127]), .B(Output1[127]), .S0(dec), .Y(n1287) );
  XNOR2X1 U5569 ( .A(n1772), .B(n4621), .Y(Output1[127]) );
  NOR2X1 U5570 ( .A(n253), .B(n4619), .Y(n4621) );
  AOI221XL U5571 ( .A0(n2152), .A1(n291), .B0(n295), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_D1[121]), .C0(n4622), .Y(n1772) );
  CLKINVX1 U5572 ( .A(n4623), .Y(n4622) );
  AOI222XL U5573 ( .A0(n2312), .A1(n4624), .B0(n2258), .B1(n4625), .C0(n264), 
        .C1(n4626), .Y(n4623) );
  XOR2X1 U5574 ( .A(n4581), .B(n4419), .Y(n4626) );
  XOR2X1 U5575 ( .A(n3630), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[40]), .Y(
        n4419) );
  XNOR2X1 U5576 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[120]), .B(n4627), .Y(
        n3630) );
  CLKINVX1 U5577 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[16]), .Y(n4581) );
  XOR2X1 U5578 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[88]), .B(n4628), .Y(
        n4625) );
  CLKINVX1 U5579 ( .A(Input1[127]), .Y(n4619) );
  CLKINVX1 U5580 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_127_), .Y(n4618) );
  OAI221X1 U5581 ( .A0(n1291), .A1(n166), .B0(n1773), .B1(n154), .C0(n4629), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_126_N3) );
  AOI22XL U5582 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_126_), 
        .B0(n221), .B1(Input1[126]), .Y(n4629) );
  MXI2X1 U5583 ( .A(Input1[126]), .B(Output1[126]), .S0(dec), .Y(n1291) );
  XOR2X1 U5584 ( .A(n4630), .B(n1773), .Y(Output1[126]) );
  CLKINVX1 U5585 ( .A(n4631), .Y(n1773) );
  OAI221X1 U5586 ( .A0(n4632), .A1(n2273), .B0(n4633), .B1(n2274), .C0(n4634), 
        .Y(n4631) );
  AOI22XL U5587 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[122]), .A1(n298), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D1[121]), .B1(n292), .Y(n4634) );
  XOR2X1 U5588 ( .A(n4635), .B(n4636), .Y(n4633) );
  MXI2X1 U5589 ( .A(n4522), .B(n4637), .S0(n314), .Y(n4636) );
  XOR2X1 U5590 ( .A(n3647), .B(n4638), .Y(n4637) );
  CLKINVX1 U5591 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[92]), .Y(n3647) );
  CLKNAND2X2 U5592 ( .A(n2148), .B(n2029), .Y(n4635) );
  XOR2X1 U5593 ( .A(n4428), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[20]), .Y(
        n4632) );
  XOR2X1 U5594 ( .A(n3643), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[44]), .Y(
        n4428) );
  XOR2X1 U5595 ( .A(n4522), .B(n4639), .Y(n3643) );
  CLKINVX1 U5596 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[124]), .Y(n4522) );
  CLKNAND2X2 U5597 ( .A(Input1[126]), .B(n2288), .Y(n4630) );
  OAI221X1 U5598 ( .A0(n1294), .A1(n166), .B0(n1774), .B1(n154), .C0(n4640), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_125_N3) );
  AOI22XL U5599 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_125_), 
        .B0(n221), .B1(Input1[125]), .Y(n4640) );
  MXI2X1 U5600 ( .A(Input1[125]), .B(Output1[125]), .S0(dec), .Y(n1294) );
  XOR2X1 U5601 ( .A(n4641), .B(n1774), .Y(Output1[125]) );
  CLKINVX1 U5602 ( .A(n4642), .Y(n1774) );
  OAI222X1 U5603 ( .A0(n4643), .A1(n2274), .B0(n4644), .B1(n2273), .C0(n2730), 
        .C1(n4645), .Y(n4642) );
  CLKINVX1 U5604 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .Y(n4645) );
  XOR2X1 U5605 ( .A(n4452), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[16]), .Y(
        n4644) );
  XOR2X1 U5606 ( .A(n3660), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[40]), .Y(
        n4452) );
  XOR2X1 U5607 ( .A(n4532), .B(n4628), .Y(n3660) );
  XOR2X1 U5608 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[53]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_53_), .Y(n4628) );
  XOR2X1 U5609 ( .A(n4646), .B(n4647), .Y(n4643) );
  MXI2X1 U5610 ( .A(n4532), .B(n4648), .S0(n314), .Y(n4647) );
  XOR2X1 U5611 ( .A(n1996), .B(n4649), .Y(n4648) );
  XOR2X1 U5612 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[88]), .B(n4650), .Y(
        n4649) );
  CLKINVX1 U5613 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[120]), .Y(n4532) );
  CLKNAND2X2 U5614 ( .A(n4651), .B(n4652), .Y(n4646) );
  CLKNAND2X2 U5615 ( .A(Input1[125]), .B(n2288), .Y(n4641) );
  OAI221X1 U5616 ( .A0(n1297), .A1(n166), .B0(n1775), .B1(n154), .C0(n4653), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_124_N3) );
  AOI22XL U5617 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_124_), 
        .B0(n221), .B1(Input1[124]), .Y(n4653) );
  MXI2X1 U5618 ( .A(Input1[124]), .B(Output1[124]), .S0(dec), .Y(n1297) );
  XNOR2X1 U5619 ( .A(n1775), .B(n4654), .Y(Output1[124]) );
  NOR2BX1 U5620 ( .AN(Input1[124]), .B(n254), .Y(n4654) );
  AOI221XL U5621 ( .A0(n2031), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .C0(n4655), .Y(n1775) );
  AO22X1 U5622 ( .A0(n268), .A1(n4656), .B0(n301), .B1(n4657), .Y(n4655) );
  XOR2X1 U5623 ( .A(n4464), .B(n2014), .Y(n4656) );
  XOR2X1 U5624 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_5_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[19]), .Y(n2014) );
  XOR2X1 U5625 ( .A(n3676), .B(n2110), .Y(n4464) );
  XOR2X1 U5626 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_11_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[43]), .Y(n2110) );
  XOR2X1 U5627 ( .A(n4638), .B(n2033), .Y(n3676) );
  XOR2X1 U5628 ( .A(n4658), .B(n4659), .Y(n4638) );
  CLKINVX1 U5629 ( .A(n4651), .Y(n2031) );
  MXI2X1 U5630 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[123]), .B(n4660), .S0(
        n314), .Y(n4651) );
  XOR2X1 U5631 ( .A(n1994), .B(n4661), .Y(n4660) );
  XOR2X1 U5632 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[91]), .B(n4662), .Y(
        n4661) );
  OAI221X1 U5633 ( .A0(n1300), .A1(n166), .B0(n4663), .B1(n154), .C0(n4664), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_123_N3) );
  AOI22XL U5634 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_123_), 
        .B0(n220), .B1(Input1[123]), .Y(n4664) );
  CLKINVX1 U5635 ( .A(n1777), .Y(n4663) );
  MXI2X1 U5636 ( .A(Input1[123]), .B(Output1[123]), .S0(dec), .Y(n1300) );
  XOR2X1 U5637 ( .A(n1777), .B(n4665), .Y(Output1[123]) );
  NOR2BX1 U5638 ( .AN(Input1[123]), .B(n255), .Y(n4665) );
  OAI2B11X1 U5639 ( .A1N(Inst_forkAE_CipherInst_RF_S_MID_D1[122]), .A0(n2255), 
        .B0(n4666), .C0(n4667), .Y(n1777) );
  AOI22XL U5640 ( .A0(n2258), .A1(n4668), .B0(n260), .B1(n4669), .Y(n4667) );
  XOR2X1 U5641 ( .A(n4508), .B(n4470), .Y(n4669) );
  XOR2X1 U5642 ( .A(n3685), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[41]), .Y(
        n4470) );
  XOR2X1 U5643 ( .A(n4670), .B(n4671), .Y(n3685) );
  XOR2X1 U5644 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[121]), .B(n4662), .Y(
        n4671) );
  XOR2X1 U5645 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[51]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_51_), .Y(n4662) );
  CLKINVX1 U5646 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[17]), .Y(n4508) );
  XOR2X1 U5647 ( .A(Inst_forkAE_CipherInst_ROUND_CST[2]), .B(n4672), .Y(n4668)
         );
  XOR2X1 U5648 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[90]), .B(n4673), .Y(
        n4672) );
  CLKINVX1 U5649 ( .A(n4674), .Y(Inst_forkAE_CipherInst_ROUND_CST[2]) );
  MXI2X1 U5650 ( .A(n4675), .B(n4676), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[124]), .Y(n4666) );
  OAI21X1 U5651 ( .A0(n4677), .A1(n283), .B0(n2267), .Y(n4676) );
  NOR2X1 U5652 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .Y(n4677) );
  NOR3X1 U5653 ( .A(n2266), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .Y(n4675) );
  OAI221X1 U5654 ( .A0(n1303), .A1(n166), .B0(n4678), .B1(n154), .C0(n4679), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_122_N3) );
  AOI22XL U5655 ( .A0(n192), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_122_), 
        .B0(n220), .B1(Input1[122]), .Y(n4679) );
  CLKINVX1 U5656 ( .A(n1779), .Y(n4678) );
  MXI2X1 U5657 ( .A(Input1[122]), .B(Output1[122]), .S0(dec), .Y(n1303) );
  XOR2X1 U5658 ( .A(n1779), .B(n4680), .Y(Output1[122]) );
  NOR2BX1 U5659 ( .AN(Input1[122]), .B(n255), .Y(n4680) );
  OAI221X1 U5660 ( .A0(n4681), .A1(n2273), .B0(n2148), .B1(n2274), .C0(n4682), 
        .Y(n1779) );
  MXI2X1 U5661 ( .A(n4683), .B(n4684), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[120]), .Y(n4682) );
  OAI21X1 U5662 ( .A0(n4685), .A1(n283), .B0(n2267), .Y(n4684) );
  NOR2X1 U5663 ( .A(n2033), .B(n2152), .Y(n4685) );
  NOR3X1 U5664 ( .A(n274), .B(n2033), .C(n2152), .Y(n4683) );
  MXI2X1 U5665 ( .A(n4657), .B(n4686), .S0(n315), .Y(n2148) );
  XOR2X1 U5666 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[92]), .B(n4639), .Y(
        n4686) );
  XOR2X1 U5667 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[54]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_54_), .Y(n4639) );
  XOR2X1 U5668 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_31_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .Y(n4657) );
  XOR2X1 U5669 ( .A(n4481), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .Y(
        n4681) );
  XOR2X1 U5670 ( .A(n3699), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[44]), .Y(
        n4481) );
  XOR2X1 U5671 ( .A(n4674), .B(n4687), .Y(n3699) );
  XOR2X1 U5672 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[124]), .B(n4673), .Y(
        n4687) );
  XOR2X1 U5673 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[50]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_50_), .Y(n4673) );
  MXI2X1 U5674 ( .A(n464), .B(n461), .S0(n1989), .Y(n4674) );
  OAI221X1 U5675 ( .A0(n1306), .A1(n179), .B0(n1780), .B1(n154), .C0(n4688), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_121_N3) );
  AOI22XL U5676 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_121_), 
        .B0(n220), .B1(Input1[121]), .Y(n4688) );
  MXI2X1 U5677 ( .A(Input1[121]), .B(Output1[121]), .S0(dec), .Y(n1306) );
  XOR2X1 U5678 ( .A(n4689), .B(n1780), .Y(Output1[121]) );
  CLKINVX1 U5679 ( .A(n4690), .Y(n1780) );
  OAI221X1 U5680 ( .A0(n2273), .A1(n4691), .B0(n2029), .B1(n2274), .C0(n4692), 
        .Y(n4690) );
  AOI22XL U5681 ( .A0(n291), .A1(n2033), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[123]), .B1(n300), .Y(n4692) );
  XOR2X1 U5682 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_31_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[123]), .Y(n2033) );
  MXI2X1 U5683 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .B(n4693), .S0(
        n315), .Y(n2029) );
  XOR2X1 U5684 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[95]), .B(n4627), .Y(
        n4693) );
  XOR2X1 U5685 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[55]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_55_), .Y(n4627) );
  XNOR2X1 U5686 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[23]), .B(n4490), .Y(
        n4691) );
  XNOR2X1 U5687 ( .A(n3718), .B(n4276), .Y(n4490) );
  CLKINVX1 U5688 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[47]), .Y(n4276) );
  XOR2X1 U5689 ( .A(n5718), .B(n4694), .Y(n3718) );
  XOR2X1 U5690 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[127]), .B(n4695), .Y(
        n4694) );
  CLKNAND2X2 U5691 ( .A(Input1[121]), .B(n2288), .Y(n4689) );
  OAI221X1 U5692 ( .A0(n1309), .A1(n171), .B0(n1781), .B1(n156), .C0(n4696), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_120_N3) );
  AOI22XL U5693 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_120_), 
        .B0(n220), .B1(Input1[120]), .Y(n4696) );
  MXI2X1 U5694 ( .A(Input1[120]), .B(Output1[120]), .S0(dec), .Y(n1309) );
  XNOR2X1 U5695 ( .A(n1781), .B(n4697), .Y(Output1[120]) );
  NOR2BX1 U5696 ( .AN(Input1[120]), .B(n255), .Y(n4697) );
  AOI221XL U5697 ( .A0(n2150), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[120]), .C0(n4698), .Y(n1781) );
  AO22X1 U5698 ( .A0(n268), .A1(n4699), .B0(n301), .B1(n4624), .Y(n4698) );
  XOR2X1 U5699 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_30_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[120]), .Y(n4624) );
  XOR2X1 U5700 ( .A(n4499), .B(n2132), .Y(n4699) );
  XOR2X1 U5701 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_4_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[18]), .Y(n2132) );
  XNOR2X1 U5702 ( .A(n3727), .B(n4251), .Y(n4499) );
  XNOR2X1 U5703 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_10_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[42]), .Y(n4251) );
  XNOR2X1 U5704 ( .A(n1996), .B(n4700), .Y(n3727) );
  XOR2X1 U5705 ( .A(n2152), .B(n4650), .Y(n4700) );
  XOR2X1 U5706 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[48]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_48_), .Y(n4650) );
  XOR2X1 U5707 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_30_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[122]), .Y(n2152) );
  CLKINVX1 U5708 ( .A(n4652), .Y(n2150) );
  MXI2X1 U5709 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[121]), .B(n4701), .S0(
        n315), .Y(n4652) );
  XOR2X1 U5710 ( .A(n5718), .B(n4702), .Y(n4701) );
  XOR2X1 U5711 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[89]), .B(n4695), .Y(
        n4702) );
  XOR2X1 U5712 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[49]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_49_), .Y(n4695) );
  MXI2X1 U5713 ( .A(n4703), .B(Inst_forkAE_CipherInst_CL_n27), .S0(n1989), .Y(
        n5718) );
  CLKINVX1 U5714 ( .A(Inst_forkAE_CipherInst_CL_STATE_0_), .Y(n4703) );
  OAI221X1 U5715 ( .A0(n1726), .A1(n172), .B0(n1948), .B1(n154), .C0(n4704), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_12_N3) );
  AOI22XL U5716 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_12_), 
        .B0(n220), .B1(Input1[12]), .Y(n4704) );
  CLKINVX1 U5717 ( .A(n1727), .Y(n1726) );
  OAI2B2X1 U5718 ( .A1N(Input1[12]), .A0(n2381), .B0(n4705), .B1(n2379), .Y(
        n1727) );
  CLKINVX1 U5719 ( .A(Output1[12]), .Y(n4705) );
  XOR2X1 U5720 ( .A(n4706), .B(n1948), .Y(Output1[12]) );
  AOI221XL U5721 ( .A0(n4707), .A1(n297), .B0(n2019), .B1(n2293), .C0(n4708), 
        .Y(n1948) );
  AO22X1 U5722 ( .A0(n267), .A1(n4709), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .B1(n292), .Y(n4708) );
  CLKINVX1 U5723 ( .A(n4616), .Y(n2019) );
  MXI2X1 U5724 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[11]), .B(n4710), .S0(
        n315), .Y(n4616) );
  XOR2X1 U5725 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[19]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[115]), .Y(n4710) );
  CLKNAND2X2 U5726 ( .A(Input1[12]), .B(n2288), .Y(n4706) );
  OAI221X1 U5727 ( .A0(n4711), .A1(n2300), .B0(n4712), .B1(n2302), .C0(n4713), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_119_N3) );
  AOI22XL U5728 ( .A0(n186), .A1(n1312), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1783), .Y(n4713) );
  CLKNAND2X2 U5729 ( .A(n4714), .B(n4715), .Y(n1312) );
  MXI2X1 U5730 ( .A(Input1[119]), .B(Output1[119]), .S0(dec), .Y(n4714) );
  XOR2X1 U5731 ( .A(n1783), .B(n4716), .Y(Output1[119]) );
  NOR2X1 U5732 ( .A(n253), .B(n4712), .Y(n4716) );
  OAI221X1 U5733 ( .A0(n4717), .A1(n277), .B0(n2267), .B1(n4718), .C0(n4719), 
        .Y(n1783) );
  AOI222XL U5734 ( .A0(n2312), .A1(n4720), .B0(n2258), .B1(n4721), .C0(n264), 
        .C1(n4722), .Y(n4719) );
  XOR2X1 U5735 ( .A(n3842), .B(n4507), .Y(n4722) );
  XOR2X1 U5736 ( .A(n3742), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[32]), .Y(
        n4507) );
  XNOR2X1 U5737 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[112]), .B(n4723), .Y(
        n3742) );
  CLKINVX1 U5738 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[8]), .Y(n3842) );
  XOR2X1 U5739 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[80]), .B(n4724), .Y(
        n4721) );
  CLKINVX1 U5740 ( .A(n2160), .Y(n4717) );
  CLKINVX1 U5741 ( .A(Input1[119]), .Y(n4712) );
  CLKINVX1 U5742 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_119_), .Y(n4711) );
  OAI221X1 U5743 ( .A0(n1315), .A1(n173), .B0(n1784), .B1(n154), .C0(n4725), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_118_N3) );
  AOI22XL U5744 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_118_), 
        .B0(n220), .B1(Input1[118]), .Y(n4725) );
  CLKINVX1 U5745 ( .A(n1316), .Y(n1315) );
  OAI2B2X1 U5746 ( .A1N(Output1[118]), .A0(n3350), .B0(n4726), .B1(n3351), .Y(
        n1316) );
  CLKINVX1 U5747 ( .A(Input1[118]), .Y(n4726) );
  XOR2X1 U5748 ( .A(n4727), .B(n1784), .Y(Output1[118]) );
  CLKINVX1 U5749 ( .A(n4728), .Y(n1784) );
  OAI221X1 U5750 ( .A0(n4729), .A1(n2273), .B0(n4730), .B1(n2274), .C0(n4731), 
        .Y(n4728) );
  AOI22XL U5751 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[114]), .A1(n299), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D1[113]), .B1(n291), .Y(n4731) );
  XOR2X1 U5752 ( .A(n4732), .B(n4733), .Y(n4730) );
  MXI2X1 U5753 ( .A(n4604), .B(n4734), .S0(n315), .Y(n4733) );
  XOR2X1 U5754 ( .A(n3759), .B(n4735), .Y(n4734) );
  CLKINVX1 U5755 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[84]), .Y(n3759) );
  CLKNAND2X2 U5756 ( .A(n2156), .B(n2037), .Y(n4732) );
  XOR2X1 U5757 ( .A(n4517), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[12]), .Y(
        n4729) );
  XOR2X1 U5758 ( .A(n3755), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[36]), .Y(
        n4517) );
  XOR2X1 U5759 ( .A(n4604), .B(n4736), .Y(n3755) );
  CLKINVX1 U5760 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[116]), .Y(n4604) );
  CLKNAND2X2 U5761 ( .A(Input1[118]), .B(n2288), .Y(n4727) );
  OAI221X1 U5762 ( .A0(n1319), .A1(n176), .B0(n1785), .B1(n153), .C0(n4737), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_117_N3) );
  AOI22XL U5763 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_117_), 
        .B0(n220), .B1(Input1[117]), .Y(n4737) );
  CLKINVX1 U5764 ( .A(n1320), .Y(n1319) );
  OAI2B2X1 U5765 ( .A1N(Output1[117]), .A0(n3350), .B0(n4738), .B1(n3351), .Y(
        n1320) );
  CLKINVX1 U5766 ( .A(Input1[117]), .Y(n4738) );
  XOR2X1 U5767 ( .A(n4739), .B(n1785), .Y(Output1[117]) );
  CLKINVX1 U5768 ( .A(n4740), .Y(n1785) );
  OAI222X1 U5769 ( .A0(n4741), .A1(n2274), .B0(n4742), .B1(n2273), .C0(n2730), 
        .C1(n4743), .Y(n4740) );
  XOR2X1 U5770 ( .A(n4528), .B(n4613), .Y(n4742) );
  CLKINVX1 U5771 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[8]), .Y(n4613) );
  XNOR2X1 U5772 ( .A(n3771), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[32]), .Y(
        n4528) );
  XOR2X1 U5773 ( .A(n4615), .B(n4724), .Y(n3771) );
  XOR2X1 U5774 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[5]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_5_), .Y(n4724) );
  XOR2X1 U5775 ( .A(n4744), .B(n4745), .Y(n4741) );
  MXI2X1 U5776 ( .A(n4615), .B(n4746), .S0(n315), .Y(n4745) );
  XOR2X1 U5777 ( .A(n3774), .B(n4747), .Y(n4746) );
  CLKINVX1 U5778 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[80]), .Y(n3774) );
  CLKINVX1 U5779 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[112]), .Y(n4615) );
  CLKNAND2X2 U5780 ( .A(n4748), .B(n4749), .Y(n4744) );
  CLKNAND2X2 U5781 ( .A(Input1[117]), .B(n2288), .Y(n4739) );
  OAI221X1 U5782 ( .A0(n1323), .A1(n174), .B0(n1786), .B1(n153), .C0(n4750), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_116_N3) );
  AOI22XL U5783 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_116_), 
        .B0(n220), .B1(Input1[116]), .Y(n4750) );
  CLKINVX1 U5784 ( .A(n1324), .Y(n1323) );
  OAI2B2X1 U5785 ( .A1N(Output1[116]), .A0(n3350), .B0(n4751), .B1(n3351), .Y(
        n1324) );
  XNOR2X1 U5786 ( .A(n1786), .B(n4752), .Y(Output1[116]) );
  NOR2X1 U5787 ( .A(n253), .B(n4751), .Y(n4752) );
  CLKINVX1 U5788 ( .A(Input1[116]), .Y(n4751) );
  AOI221XL U5789 ( .A0(n2039), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .C0(n4753), .Y(n1786) );
  AO22X1 U5790 ( .A0(n268), .A1(n4754), .B0(n301), .B1(n4755), .Y(n4753) );
  XOR2X1 U5791 ( .A(n2021), .B(n4540), .Y(n4754) );
  XOR2X1 U5792 ( .A(n3786), .B(n2117), .Y(n4540) );
  XOR2X1 U5793 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_9_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[35]), .Y(n2117) );
  XOR2X1 U5794 ( .A(n4735), .B(n2041), .Y(n3786) );
  XOR2X1 U5795 ( .A(n4756), .B(n4757), .Y(n4735) );
  CLKINVX1 U5796 ( .A(n4748), .Y(n2039) );
  MXI2X1 U5797 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[115]), .B(n4758), .S0(
        n315), .Y(n4748) );
  XOR2X1 U5798 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[83]), .B(n4759), .Y(
        n4758) );
  OAI221X1 U5799 ( .A0(n1327), .A1(n175), .B0(n4760), .B1(n153), .C0(n4761), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_115_N3) );
  AOI22XL U5800 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_115_), 
        .B0(n220), .B1(Input1[115]), .Y(n4761) );
  CLKINVX1 U5801 ( .A(n1788), .Y(n4760) );
  CLKINVX1 U5802 ( .A(n1328), .Y(n1327) );
  OAI2B2X1 U5803 ( .A1N(Output1[115]), .A0(n3350), .B0(n4762), .B1(n3351), .Y(
        n1328) );
  XOR2X1 U5804 ( .A(n1788), .B(n4763), .Y(Output1[115]) );
  NOR2X1 U5805 ( .A(n253), .B(n4762), .Y(n4763) );
  CLKINVX1 U5806 ( .A(Input1[115]), .Y(n4762) );
  OAI2B11X1 U5807 ( .A1N(Inst_forkAE_CipherInst_RF_S_MID_D1[114]), .A0(n2255), 
        .B0(n4764), .C0(n4765), .Y(n1788) );
  AOI22XL U5808 ( .A0(n2258), .A1(n4766), .B0(n261), .B1(n4767), .Y(n4765) );
  XOR2X1 U5809 ( .A(n4148), .B(n4554), .Y(n4767) );
  XOR2X1 U5810 ( .A(n3795), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[33]), .Y(
        n4554) );
  XOR2X1 U5811 ( .A(n4718), .B(n4759), .Y(n3795) );
  XOR2X1 U5812 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[3]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_3_), .Y(n4759) );
  CLKINVX1 U5813 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[113]), .Y(n4718) );
  CLKINVX1 U5814 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[9]), .Y(n4148) );
  XOR2X1 U5815 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[82]), .B(n4768), .Y(
        n4766) );
  MXI2X1 U5816 ( .A(n4769), .B(n4770), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[116]), .Y(n4764) );
  OAI21X1 U5817 ( .A0(n4771), .A1(n282), .B0(n2267), .Y(n4770) );
  NOR2X1 U5818 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .Y(n4771) );
  NOR3X1 U5819 ( .A(n2266), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .Y(n4769) );
  OAI221X1 U5820 ( .A0(n1331), .A1(n168), .B0(n4772), .B1(n153), .C0(n4773), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_114_N3) );
  AOI22XL U5821 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_114_), 
        .B0(n220), .B1(Input1[114]), .Y(n4773) );
  CLKINVX1 U5822 ( .A(n1790), .Y(n4772) );
  CLKINVX1 U5823 ( .A(n1332), .Y(n1331) );
  OAI2B2X1 U5824 ( .A1N(Output1[114]), .A0(n3350), .B0(n4774), .B1(n3351), .Y(
        n1332) );
  XOR2X1 U5825 ( .A(n1790), .B(n4775), .Y(Output1[114]) );
  NOR2X1 U5826 ( .A(n253), .B(n4774), .Y(n4775) );
  CLKINVX1 U5827 ( .A(Input1[114]), .Y(n4774) );
  OAI221X1 U5828 ( .A0(n4776), .A1(n2273), .B0(n2156), .B1(n2274), .C0(n4777), 
        .Y(n1790) );
  MXI2X1 U5829 ( .A(n4778), .B(n4779), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[112]), .Y(n4777) );
  OAI21X1 U5830 ( .A0(n4780), .A1(n283), .B0(n2267), .Y(n4779) );
  NOR2X1 U5831 ( .A(n2041), .B(n2160), .Y(n4780) );
  NOR3X1 U5832 ( .A(n2266), .B(n2041), .C(n2160), .Y(n4778) );
  MXI2X1 U5833 ( .A(n4755), .B(n4781), .S0(n315), .Y(n2156) );
  XOR2X1 U5834 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[84]), .B(n4736), .Y(
        n4781) );
  XOR2X1 U5835 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[6]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_6_), .Y(n4736) );
  XOR2X1 U5836 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_29_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .Y(n4755) );
  XOR2X1 U5837 ( .A(n4565), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .Y(
        n4776) );
  XOR2X1 U5838 ( .A(n3809), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[36]), .Y(
        n4565) );
  XNOR2X1 U5839 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .B(n4768), .Y(
        n3809) );
  XOR2X1 U5840 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[2]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_2_), .Y(n4768) );
  OAI221X1 U5841 ( .A0(n1335), .A1(n169), .B0(n1791), .B1(n153), .C0(n4782), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_113_N3) );
  AOI22XL U5842 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_113_), 
        .B0(n220), .B1(Input1[113]), .Y(n4782) );
  CLKINVX1 U5843 ( .A(n1336), .Y(n1335) );
  OAI2B2X1 U5844 ( .A1N(Output1[113]), .A0(n3350), .B0(n4783), .B1(n3351), .Y(
        n1336) );
  CLKINVX1 U5845 ( .A(Input1[113]), .Y(n4783) );
  XOR2X1 U5846 ( .A(n4784), .B(n1791), .Y(Output1[113]) );
  CLKINVX1 U5847 ( .A(n4785), .Y(n1791) );
  OAI221X1 U5848 ( .A0(n4786), .A1(n2273), .B0(n2037), .B1(n2274), .C0(n4787), 
        .Y(n4785) );
  AOI22XL U5849 ( .A0(n291), .A1(n2041), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[115]), .B1(n300), .Y(n4787) );
  XOR2X1 U5850 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_29_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[115]), .Y(n2041) );
  MXI2X1 U5851 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .B(n4788), .S0(
        n315), .Y(n2037) );
  XOR2X1 U5852 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[87]), .B(n4723), .Y(
        n4788) );
  XOR2X1 U5853 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[7]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_7_), .Y(n4723) );
  XNOR2X1 U5854 ( .A(n4575), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .Y(
        n4786) );
  XOR2X1 U5855 ( .A(n3822), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[39]), .Y(
        n4575) );
  XNOR2X1 U5856 ( .A(n4743), .B(n4789), .Y(n3822) );
  CLKINVX1 U5857 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[119]), .Y(n4743) );
  CLKNAND2X2 U5858 ( .A(Input1[113]), .B(n2288), .Y(n4784) );
  OAI221X1 U5859 ( .A0(n1339), .A1(n170), .B0(n1792), .B1(n153), .C0(n4790), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_112_N3) );
  AOI22XL U5860 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_112_), 
        .B0(n220), .B1(Input1[112]), .Y(n4790) );
  CLKINVX1 U5861 ( .A(n1340), .Y(n1339) );
  OAI2B2X1 U5862 ( .A1N(Output1[112]), .A0(n3350), .B0(n4791), .B1(n3351), .Y(
        n1340) );
  CLKNAND2X2 U5863 ( .A(n4715), .B(n3734), .Y(n3351) );
  CLKNAND2X2 U5864 ( .A(dec), .B(n4715), .Y(n3350) );
  CLKNAND2X2 U5865 ( .A(n4792), .B(n4238), .Y(n4715) );
  XNOR2X1 U5866 ( .A(n1792), .B(n4793), .Y(Output1[112]) );
  NOR2X1 U5867 ( .A(n253), .B(n4791), .Y(n4793) );
  CLKINVX1 U5868 ( .A(Input1[112]), .Y(n4791) );
  AOI221XL U5869 ( .A0(n2158), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[112]), .C0(n4794), .Y(n1792) );
  AO22X1 U5870 ( .A0(n268), .A1(n4795), .B0(n301), .B1(n4720), .Y(n4794) );
  XOR2X1 U5871 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_28_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[112]), .Y(n4720) );
  XOR2X1 U5872 ( .A(n4582), .B(n2140), .Y(n4795) );
  XNOR2X1 U5873 ( .A(n3831), .B(n4339), .Y(n4582) );
  XNOR2X1 U5874 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_8_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[34]), .Y(n4339) );
  XOR2X1 U5875 ( .A(n4747), .B(n2160), .Y(n3831) );
  XOR2X1 U5876 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_28_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[114]), .Y(n2160) );
  XOR2X1 U5877 ( .A(n4796), .B(n4797), .Y(n4747) );
  CLKINVX1 U5878 ( .A(n4749), .Y(n2158) );
  MXI2X1 U5879 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[113]), .B(n4798), .S0(
        n315), .Y(n4749) );
  XOR2X1 U5880 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[81]), .B(n4789), .Y(
        n4798) );
  XOR2X1 U5881 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[1]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_1_), .Y(n4789) );
  OAI221X1 U5882 ( .A0(n4799), .A1(n2300), .B0(n4800), .B1(n2302), .C0(n4801), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_111_N3) );
  AOI22XL U5883 ( .A0(n186), .A1(n1343), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1794), .Y(n4801) );
  OAI222X1 U5884 ( .A0(n4800), .A1(n3433), .B0(n3432), .B1(n4802), .C0(n4238), 
        .C1(n4803), .Y(n1343) );
  CLKINVX1 U5885 ( .A(Output1[111]), .Y(n4802) );
  XOR2X1 U5886 ( .A(n1794), .B(n4804), .Y(Output1[111]) );
  NOR2X1 U5887 ( .A(n254), .B(n4800), .Y(n4804) );
  OAI221X1 U5888 ( .A0(n4805), .A1(n277), .B0(n2267), .B1(n4806), .C0(n4807), 
        .Y(n1794) );
  AOI222XL U5889 ( .A0(n2312), .A1(n4808), .B0(n2258), .B1(n4809), .C0(n264), 
        .C1(n4810), .Y(n4807) );
  XOR2X1 U5890 ( .A(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]), .B(n4592), .Y(
        n4810) );
  XNOR2X1 U5891 ( .A(n3851), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[56]), .Y(
        n4592) );
  XNOR2X1 U5892 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[104]), .B(n4811), .Y(
        n3851) );
  XOR2X1 U5893 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[72]), .B(n4812), .Y(
        n4809) );
  CLKINVX1 U5894 ( .A(n2172), .Y(n4805) );
  CLKINVX1 U5895 ( .A(Input1[111]), .Y(n4800) );
  CLKINVX1 U5896 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_111_), .Y(n4799) );
  OAI221X1 U5897 ( .A0(n1346), .A1(n165), .B0(n1795), .B1(n153), .C0(n4813), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_110_N3) );
  AOI22XL U5898 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_110_), 
        .B0(n220), .B1(Input1[110]), .Y(n4813) );
  CLKINVX1 U5899 ( .A(n1347), .Y(n1346) );
  OAI2B2X1 U5900 ( .A1N(Output1[110]), .A0(n3432), .B0(n4814), .B1(n3433), .Y(
        n1347) );
  CLKINVX1 U5901 ( .A(Input1[110]), .Y(n4814) );
  XOR2X1 U5902 ( .A(n4815), .B(n1795), .Y(Output1[110]) );
  CLKINVX1 U5903 ( .A(n4816), .Y(n1795) );
  OAI221X1 U5904 ( .A0(n4817), .A1(n2273), .B0(n4818), .B1(n2274), .C0(n4819), 
        .Y(n4816) );
  AOI22XL U5905 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[106]), .A1(n299), 
        .B0(Inst_forkAE_CipherInst_RF_S_MID_D1[105]), .B1(n292), .Y(n4819) );
  XOR2X1 U5906 ( .A(n4820), .B(n4821), .Y(n4818) );
  MXI2X1 U5907 ( .A(n4112), .B(n4822), .S0(n315), .Y(n4821) );
  XOR2X1 U5908 ( .A(n3868), .B(n4823), .Y(n4822) );
  CLKINVX1 U5909 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[76]), .Y(n3868) );
  CLKNAND2X2 U5910 ( .A(n2164), .B(n2045), .Y(n4820) );
  XOR2X1 U5911 ( .A(n4599), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[4]), .Y(
        n4817) );
  XOR2X1 U5912 ( .A(n3864), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[60]), .Y(
        n4599) );
  XOR2X1 U5913 ( .A(n4112), .B(n4824), .Y(n3864) );
  CLKINVX1 U5914 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[108]), .Y(n4112) );
  CLKNAND2X2 U5915 ( .A(Input1[110]), .B(n2288), .Y(n4815) );
  OAI221X1 U5916 ( .A0(n1730), .A1(n167), .B0(n4825), .B1(n153), .C0(n4826), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_11_N3) );
  AOI22XL U5917 ( .A0(n191), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_11_), 
        .B0(n219), .B1(Input1[11]), .Y(n4826) );
  CLKINVX1 U5918 ( .A(n1950), .Y(n4825) );
  CLKINVX1 U5919 ( .A(n1731), .Y(n1730) );
  OAI2B2X1 U5920 ( .A1N(Output1[11]), .A0(n2379), .B0(n4827), .B1(n2381), .Y(
        n1731) );
  XOR2X1 U5921 ( .A(n1950), .B(n4828), .Y(Output1[11]) );
  NOR2X1 U5922 ( .A(n253), .B(n4827), .Y(n4828) );
  CLKINVX1 U5923 ( .A(Input1[11]), .Y(n4827) );
  OAI211XL U5924 ( .A0(n4829), .A1(n2273), .B0(n4830), .C0(n4831), .Y(n1950)
         );
  AOI22XL U5925 ( .A0(n2258), .A1(n4832), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[10]), .B1(n2312), .Y(n4831) );
  XOR2X1 U5926 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[18]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[114]), .Y(n4832) );
  MXI2X1 U5927 ( .A(n4833), .B(n4834), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[12]), .Y(n4830) );
  OAI21X1 U5928 ( .A0(n4835), .A1(n283), .B0(n2267), .Y(n4834) );
  NOR2X1 U5929 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .Y(n4835) );
  NOR3X1 U5930 ( .A(n2266), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .Y(n4833) );
  OAI221X1 U5931 ( .A0(n1350), .A1(n165), .B0(n1796), .B1(n153), .C0(n4836), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_109_N3) );
  AOI22XL U5932 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_109_), 
        .B0(n219), .B1(Input1[109]), .Y(n4836) );
  CLKINVX1 U5933 ( .A(n1351), .Y(n1350) );
  OAI2B2X1 U5934 ( .A1N(Output1[109]), .A0(n3432), .B0(n4837), .B1(n3433), .Y(
        n1351) );
  CLKINVX1 U5935 ( .A(Input1[109]), .Y(n4837) );
  XOR2X1 U5936 ( .A(n4838), .B(n1796), .Y(Output1[109]) );
  CLKINVX1 U5937 ( .A(n4839), .Y(n1796) );
  OAI222X1 U5938 ( .A0(n4840), .A1(n2274), .B0(n4841), .B1(n2273), .C0(n2730), 
        .C1(n4842), .Y(n4839) );
  XOR2X1 U5939 ( .A(n4610), .B(n4185), .Y(n4841) );
  CLKINVX1 U5940 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[0]), .Y(n4185) );
  XNOR2X1 U5941 ( .A(n3880), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[56]), .Y(
        n4610) );
  XOR2X1 U5942 ( .A(n4224), .B(n4812), .Y(n3880) );
  XOR2X1 U5943 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[61]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_61_), .Y(n4812) );
  XOR2X1 U5944 ( .A(n4843), .B(n4844), .Y(n4840) );
  MXI2X1 U5945 ( .A(n4224), .B(n4845), .S0(n315), .Y(n4844) );
  XOR2X1 U5946 ( .A(n3883), .B(n4846), .Y(n4845) );
  CLKINVX1 U5947 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[72]), .Y(n3883) );
  CLKINVX1 U5948 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[104]), .Y(n4224) );
  CLKNAND2X2 U5949 ( .A(n4847), .B(n4848), .Y(n4843) );
  CLKNAND2X2 U5950 ( .A(Input1[109]), .B(n2288), .Y(n4838) );
  OAI221X1 U5951 ( .A0(n1354), .A1(n165), .B0(n1797), .B1(n153), .C0(n4849), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_108_N3) );
  AOI22XL U5952 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_108_), 
        .B0(n219), .B1(Input1[108]), .Y(n4849) );
  CLKINVX1 U5953 ( .A(n1355), .Y(n1354) );
  OAI2B2X1 U5954 ( .A1N(Output1[108]), .A0(n3432), .B0(n4850), .B1(n3433), .Y(
        n1355) );
  XNOR2X1 U5955 ( .A(n1797), .B(n4851), .Y(Output1[108]) );
  NOR2X1 U5956 ( .A(n254), .B(n4850), .Y(n4851) );
  CLKINVX1 U5957 ( .A(Input1[108]), .Y(n4850) );
  AOI221XL U5958 ( .A0(n2051), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .C0(n4852), .Y(n1797) );
  AO22X1 U5959 ( .A0(n268), .A1(n4853), .B0(n301), .B1(n4854), .Y(n4852) );
  XOR2X1 U5960 ( .A(n2049), .B(n4709), .Y(n4853) );
  XOR2X1 U5961 ( .A(n3895), .B(n2096), .Y(n4709) );
  XOR2X1 U5962 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_15_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[59]), .Y(n2096) );
  XOR2X1 U5963 ( .A(n4823), .B(n2053), .Y(n3895) );
  XOR2X1 U5964 ( .A(n4855), .B(n4856), .Y(n4823) );
  CLKINVX1 U5965 ( .A(n4847), .Y(n2051) );
  MXI2X1 U5966 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[107]), .B(n4857), .S0(
        n316), .Y(n4847) );
  XOR2X1 U5967 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[75]), .B(n4858), .Y(
        n4857) );
  OAI221X1 U5968 ( .A0(n1358), .A1(n165), .B0(n4859), .B1(n153), .C0(n4860), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_107_N3) );
  AOI22XL U5969 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_107_), 
        .B0(n219), .B1(Input1[107]), .Y(n4860) );
  CLKINVX1 U5970 ( .A(n1799), .Y(n4859) );
  CLKINVX1 U5971 ( .A(n1359), .Y(n1358) );
  OAI2B2X1 U5972 ( .A1N(Output1[107]), .A0(n3432), .B0(n4861), .B1(n3433), .Y(
        n1359) );
  XOR2X1 U5973 ( .A(n1799), .B(n4862), .Y(Output1[107]) );
  NOR2X1 U5974 ( .A(n254), .B(n4861), .Y(n4862) );
  CLKINVX1 U5975 ( .A(Input1[107]), .Y(n4861) );
  OAI2B11X1 U5976 ( .A1N(Inst_forkAE_CipherInst_RF_S_MID_D1[106]), .A0(n2255), 
        .B0(n4863), .C0(n4864), .Y(n1799) );
  AOI22XL U5977 ( .A0(n2258), .A1(n4865), .B0(n260), .B1(n4866), .Y(n4864) );
  XOR2X1 U5978 ( .A(n3980), .B(n4829), .Y(n4866) );
  XOR2X1 U5979 ( .A(n3904), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[57]), .Y(
        n4829) );
  XOR2X1 U5980 ( .A(n4806), .B(n4858), .Y(n3904) );
  XOR2X1 U5981 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[59]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_59_), .Y(n4858) );
  CLKINVX1 U5982 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[105]), .Y(n4806) );
  CLKINVX1 U5983 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[1]), .Y(n3980) );
  XOR2X1 U5984 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[74]), .B(n4867), .Y(
        n4865) );
  MXI2X1 U5985 ( .A(n4868), .B(n4869), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[108]), .Y(n4863) );
  OAI21X1 U5986 ( .A0(n4870), .A1(n283), .B0(n2267), .Y(n4869) );
  NOR2X1 U5987 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .Y(n4870) );
  NOR3X1 U5988 ( .A(n284), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .C(
        Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .Y(n4868) );
  OAI221X1 U5989 ( .A0(n1362), .A1(n165), .B0(n4871), .B1(n153), .C0(n4872), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_106_N3) );
  AOI22XL U5990 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_106_), 
        .B0(n219), .B1(Input1[106]), .Y(n4872) );
  CLKINVX1 U5991 ( .A(n1801), .Y(n4871) );
  CLKINVX1 U5992 ( .A(n1363), .Y(n1362) );
  OAI2B2X1 U5993 ( .A1N(Output1[106]), .A0(n3432), .B0(n4873), .B1(n3433), .Y(
        n1363) );
  XOR2X1 U5994 ( .A(n1801), .B(n4874), .Y(Output1[106]) );
  NOR2X1 U5995 ( .A(n253), .B(n4873), .Y(n4874) );
  CLKINVX1 U5996 ( .A(Input1[106]), .Y(n4873) );
  OAI221X1 U5997 ( .A0(n4875), .A1(n2273), .B0(n2164), .B1(n2274), .C0(n4876), 
        .Y(n1801) );
  MXI2X1 U5998 ( .A(n4877), .B(n4878), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[104]), .Y(n4876) );
  OAI21X1 U5999 ( .A0(n4879), .A1(n282), .B0(n2267), .Y(n4878) );
  NOR2X1 U6000 ( .A(n2172), .B(n2053), .Y(n4879) );
  NOR3X1 U6001 ( .A(n2266), .B(n2172), .C(n2053), .Y(n4877) );
  MXI2X1 U6002 ( .A(n4854), .B(n4880), .S0(n316), .Y(n2164) );
  XOR2X1 U6003 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[76]), .B(n4824), .Y(
        n4880) );
  XOR2X1 U6004 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[62]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_62_), .Y(n4824) );
  XOR2X1 U6005 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_27_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .Y(n4854) );
  XOR2X1 U6006 ( .A(n4881), .B(Inst_forkAE_CipherInst_RF_SHIFT1_OUT[10]), .Y(
        n4875) );
  OAI221X1 U6007 ( .A0(n1366), .A1(n165), .B0(n1802), .B1(n153), .C0(n4882), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_105_N3) );
  AOI22XL U6008 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_105_), 
        .B0(n219), .B1(Input1[105]), .Y(n4882) );
  CLKINVX1 U6009 ( .A(n1367), .Y(n1366) );
  OAI2B2X1 U6010 ( .A1N(Output1[105]), .A0(n3432), .B0(n4883), .B1(n3433), .Y(
        n1367) );
  CLKINVX1 U6011 ( .A(Input1[105]), .Y(n4883) );
  XOR2X1 U6012 ( .A(n4884), .B(n1802), .Y(Output1[105]) );
  CLKINVX1 U6013 ( .A(n4885), .Y(n1802) );
  OAI221X1 U6014 ( .A0(n2273), .A1(n4886), .B0(n2045), .B1(n2274), .C0(n4887), 
        .Y(n4885) );
  AOI22XL U6015 ( .A0(n291), .A1(n2053), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[107]), .B1(n300), .Y(n4887) );
  XOR2X1 U6016 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_27_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[107]), .Y(n2053) );
  MXI2X1 U6017 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .B(n4888), .S0(
        n316), .Y(n2045) );
  XOR2X1 U6018 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[79]), .B(n4811), .Y(
        n4888) );
  XOR2X1 U6019 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[63]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_63_), .Y(n4811) );
  XOR2X1 U6020 ( .A(n4218), .B(n3711), .Y(n4886) );
  XOR2X1 U6021 ( .A(n3931), .B(n4089), .Y(n3711) );
  CLKINVX1 U6022 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[63]), .Y(n4089) );
  XNOR2X1 U6023 ( .A(n4842), .B(n4889), .Y(n3931) );
  CLKINVX1 U6024 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .Y(n4842) );
  CLKINVX1 U6025 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .Y(n4218) );
  CLKNAND2X2 U6026 ( .A(Input1[105]), .B(n2288), .Y(n4884) );
  OAI221X1 U6027 ( .A0(n1370), .A1(n165), .B0(n1803), .B1(n153), .C0(n4890), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_104_N3) );
  AOI22XL U6028 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_104_), 
        .B0(n219), .B1(Input1[104]), .Y(n4890) );
  CLKINVX1 U6029 ( .A(n1371), .Y(n1370) );
  OAI2B2X1 U6030 ( .A1N(Output1[104]), .A0(n3432), .B0(n4891), .B1(n3433), .Y(
        n1371) );
  CLKNAND2X2 U6031 ( .A(n4803), .B(n3734), .Y(n3433) );
  CLKNAND2X2 U6032 ( .A(dec), .B(n4803), .Y(n3432) );
  XNOR2X1 U6033 ( .A(n1803), .B(n4892), .Y(Output1[104]) );
  NOR2X1 U6034 ( .A(n254), .B(n4891), .Y(n4892) );
  CLKINVX1 U6035 ( .A(Input1[104]), .Y(n4891) );
  AOI221XL U6036 ( .A0(n2170), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[104]), .C0(n4893), .Y(n1803) );
  AO22X1 U6037 ( .A0(n267), .A1(n4894), .B0(n301), .B1(n4808), .Y(n4893) );
  XOR2X1 U6038 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_26_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[104]), .Y(n4808) );
  XOR2X1 U6039 ( .A(n3843), .B(n2168), .Y(n4894) );
  XOR2X1 U6040 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_0_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[2]), .Y(n2168) );
  XOR2X1 U6041 ( .A(n3940), .B(n2219), .Y(n3843) );
  CLKINVX1 U6042 ( .A(n4064), .Y(n2219) );
  XNOR2X1 U6043 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_14_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[58]), .Y(n4064) );
  XOR2X1 U6044 ( .A(n4846), .B(n2172), .Y(n3940) );
  XOR2X1 U6045 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_26_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[106]), .Y(n2172) );
  XOR2X1 U6046 ( .A(n4895), .B(n4896), .Y(n4846) );
  CLKINVX1 U6047 ( .A(n4848), .Y(n2170) );
  MXI2X1 U6048 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[105]), .B(n4897), .S0(
        n316), .Y(n4848) );
  XOR2X1 U6049 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[73]), .B(n4889), .Y(
        n4897) );
  XOR2X1 U6050 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[57]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_57_), .Y(n4889) );
  OAI221X1 U6051 ( .A0(n4898), .A1(n2300), .B0(n4899), .B1(n2302), .C0(n4900), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_103_N3) );
  AOI22XL U6052 ( .A0(n184), .A1(n1374), .B0(
        Inst_forkAE_ControlInst_fsm_state_1_), .B1(n1805), .Y(n4900) );
  OAI222X1 U6053 ( .A0(n2250), .A1(n4901), .B0(n4902), .B1(n3949), .C0(n4899), 
        .C1(n2252), .Y(n1374) );
  CLKNAND2X2 U6054 ( .A(Block_Size[1]), .B(n4238), .Y(n3949) );
  CLKINVX1 U6055 ( .A(Output1[103]), .Y(n4901) );
  XOR2X1 U6056 ( .A(n1805), .B(n4903), .Y(Output1[103]) );
  NOR2X1 U6057 ( .A(n254), .B(n4899), .Y(n4903) );
  OAI221X1 U6058 ( .A0(n2267), .A1(n4444), .B0(n3606), .B1(n279), .C0(n4904), 
        .Y(n1805) );
  AOI222XL U6059 ( .A0(n2312), .A1(n3620), .B0(n2258), .B1(n4905), .C0(n264), 
        .C1(n4906), .Y(n4904) );
  XOR2X1 U6060 ( .A(n4498), .B(n3979), .Y(n4906) );
  XOR2X1 U6061 ( .A(n3951), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[48]), .Y(
        n3979) );
  XNOR2X1 U6062 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[96]), .B(n4907), .Y(
        n3951) );
  CLKINVX1 U6063 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[24]), .Y(n4498) );
  XOR2X1 U6064 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[64]), .B(n4908), .Y(
        n4905) );
  XOR2X1 U6065 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_24_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[96]), .Y(n3620) );
  CLKNAND2X2 U6066 ( .A(n2293), .B(n322), .Y(n2255) );
  CLKINVX1 U6067 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[97]), .Y(n4444) );
  CLKINVX1 U6068 ( .A(Input1[103]), .Y(n4899) );
  CLKINVX1 U6069 ( .A(Inst_forkAE_MainPart1_Tag_Reg_Output_103_), .Y(n4898) );
  OAI221X1 U6070 ( .A0(n1377), .A1(n165), .B0(n1806), .B1(n153), .C0(n4909), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_102_N3) );
  AOI22XL U6071 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_102_), 
        .B0(n219), .B1(Input1[102]), .Y(n4909) );
  CLKINVX1 U6072 ( .A(n1378), .Y(n1377) );
  OAI2B2X1 U6073 ( .A1N(Output1[102]), .A0(n2250), .B0(n4910), .B1(n2252), .Y(
        n1378) );
  CLKINVX1 U6074 ( .A(Input1[102]), .Y(n4910) );
  XOR2X1 U6075 ( .A(n4911), .B(n1806), .Y(Output1[102]) );
  CLKINVX1 U6076 ( .A(n4912), .Y(n1806) );
  OAI221X1 U6077 ( .A0(n4913), .A1(n2273), .B0(n4914), .B1(n2274), .C0(n4915), 
        .Y(n4912) );
  AOI22XL U6078 ( .A0(Inst_forkAE_CipherInst_RF_S_MID_D1[98]), .A1(n299), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[97]), .B1(n292), .Y(n4915) );
  XOR2X1 U6079 ( .A(n4916), .B(n4917), .Y(n4914) );
  MXI2X1 U6080 ( .A(n4433), .B(n4918), .S0(n316), .Y(n4917) );
  XOR2X1 U6081 ( .A(n3968), .B(n4919), .Y(n4918) );
  CLKINVX1 U6082 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[68]), .Y(n3968) );
  CLKNAND2X2 U6083 ( .A(n2176), .B(n2057), .Y(n4916) );
  MXI2X1 U6084 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .B(n4920), .S0(
        n316), .Y(n2057) );
  XOR2X1 U6085 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[71]), .B(n4907), .Y(
        n4920) );
  XOR2X1 U6086 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[23]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_23_), .Y(n4907) );
  MXI2X1 U6087 ( .A(n4921), .B(n4922), .S0(n316), .Y(n2176) );
  XOR2X1 U6088 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[68]), .B(n4923), .Y(
        n4922) );
  XOR2X1 U6089 ( .A(n4106), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[28]), .Y(
        n4913) );
  XOR2X1 U6090 ( .A(n3964), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[52]), .Y(
        n4106) );
  XOR2X1 U6091 ( .A(n4433), .B(n4923), .Y(n3964) );
  XOR2X1 U6092 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[22]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_22_), .Y(n4923) );
  CLKINVX1 U6093 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[100]), .Y(n4433) );
  CLKNAND2X2 U6094 ( .A(Input1[102]), .B(n2288), .Y(n4911) );
  OAI221X1 U6095 ( .A0(n1381), .A1(n165), .B0(n1807), .B1(n153), .C0(n4924), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_101_N3) );
  AOI22XL U6096 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_101_), 
        .B0(n219), .B1(Input1[101]), .Y(n4924) );
  CLKINVX1 U6097 ( .A(n1382), .Y(n1381) );
  OAI2B2X1 U6098 ( .A1N(Input1[101]), .A0(n2252), .B0(n4925), .B1(n2250), .Y(
        n1382) );
  CLKINVX1 U6099 ( .A(Output1[101]), .Y(n4925) );
  XOR2X1 U6100 ( .A(n4926), .B(n1807), .Y(Output1[101]) );
  AOI222XL U6101 ( .A0(n4927), .A1(n2293), .B0(n4928), .B1(n265), .C0(n2332), 
        .C1(Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .Y(n1807) );
  CLKINVX1 U6102 ( .A(n2730), .Y(n2332) );
  NOR2X1 U6103 ( .A(n286), .B(n294), .Y(n2730) );
  XOR2X1 U6104 ( .A(n4220), .B(n4281), .Y(n4928) );
  CLKINVX1 U6105 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[24]), .Y(n4281) );
  XOR2X1 U6106 ( .A(n3990), .B(Inst_forkAE_CipherInst_RF_S_MID_D1[48]), .Y(
        n4220) );
  XOR2X1 U6107 ( .A(n4929), .B(n4908), .Y(n3990) );
  XOR2X1 U6108 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[21]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_21_), .Y(n4908) );
  XNOR2X1 U6109 ( .A(n4930), .B(n4931), .Y(n4927) );
  MXI2X1 U6110 ( .A(n4929), .B(n4932), .S0(n316), .Y(n4931) );
  XOR2X1 U6111 ( .A(n3993), .B(n4933), .Y(n4932) );
  CLKINVX1 U6112 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[64]), .Y(n3993) );
  CLKINVX1 U6113 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[96]), .Y(n4929) );
  CLKNAND2X2 U6114 ( .A(n3622), .B(n4934), .Y(n4930) );
  MXI2X1 U6115 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[97]), .B(n4935), .S0(
        n316), .Y(n3622) );
  XOR2X1 U6116 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[65]), .B(n4936), .Y(
        n4935) );
  CLKNAND2X2 U6117 ( .A(Input1[101]), .B(n2288), .Y(n4926) );
  OAI221X1 U6118 ( .A0(n1385), .A1(n165), .B0(n1808), .B1(n152), .C0(n4937), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_100_N3) );
  AOI22XL U6119 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_100_), 
        .B0(n219), .B1(Input1[100]), .Y(n4937) );
  CLKINVX1 U6120 ( .A(n1386), .Y(n1385) );
  OAI2B2X1 U6121 ( .A1N(Output1[100]), .A0(n2250), .B0(n4938), .B1(n2252), .Y(
        n1386) );
  CLKNAND2X2 U6122 ( .A(n4902), .B(n3734), .Y(n2252) );
  CLKNAND2X2 U6123 ( .A(n4902), .B(dec), .Y(n2250) );
  AOI21X1 U6124 ( .A0(n4238), .A1(n4058), .B0(n4792), .Y(n4902) );
  CLKINVX1 U6125 ( .A(n4803), .Y(n4792) );
  CLKNAND2X2 U6126 ( .A(n4058), .B(n4057), .Y(n4803) );
  CLKINVX1 U6127 ( .A(Block_Size[1]), .Y(n4057) );
  CLKINVX1 U6128 ( .A(n3627), .Y(n4058) );
  CLKNAND2X2 U6129 ( .A(n4056), .B(n4239), .Y(n3627) );
  CLKINVX1 U6130 ( .A(Block_Size[2]), .Y(n4239) );
  CLKINVX1 U6131 ( .A(Block_Size[3]), .Y(n4056) );
  CLKINVX1 U6132 ( .A(Block_Size[0]), .Y(n4238) );
  XNOR2X1 U6133 ( .A(n1808), .B(n4939), .Y(Output1[100]) );
  NOR2X1 U6134 ( .A(n253), .B(n4938), .Y(n4939) );
  CLKINVX1 U6135 ( .A(Input1[100]), .Y(n4938) );
  AOI221XL U6136 ( .A0(n2059), .A1(n2293), .B0(n291), .B1(
        Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .C0(n4940), .Y(n1808) );
  AO22X1 U6137 ( .A0(n266), .A1(n4941), .B0(n301), .B1(n4921), .Y(n4940) );
  XOR2X1 U6138 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_25_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[100]), .Y(n4921) );
  XOR2X1 U6139 ( .A(n4332), .B(n2007), .Y(n4941) );
  XOR2X1 U6140 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_7_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[27]), .Y(n2007) );
  XOR2X1 U6141 ( .A(n2103), .B(n4005), .Y(n4332) );
  XOR2X1 U6142 ( .A(n4919), .B(n2061), .Y(n4005) );
  XOR2X1 U6143 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_25_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[99]), .Y(n2061) );
  XOR2X1 U6144 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[20]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_20_), .Y(n4919) );
  XOR2X1 U6145 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_13_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[51]), .Y(n2103) );
  CLKINVX1 U6146 ( .A(n4934), .Y(n2059) );
  MXI2X1 U6147 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[99]), .B(n4942), .S0(
        n316), .Y(n4934) );
  XOR2X1 U6148 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[67]), .B(n4445), .Y(
        n4942) );
  XOR2X1 U6149 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[19]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_19_), .Y(n4445) );
  OAI221X1 U6150 ( .A0(n1734), .A1(n165), .B0(n4943), .B1(n152), .C0(n4944), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_10_N3) );
  AOI22XL U6151 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_10_), 
        .B0(n219), .B1(Input1[10]), .Y(n4944) );
  CLKINVX1 U6152 ( .A(n1952), .Y(n4943) );
  CLKINVX1 U6153 ( .A(n1735), .Y(n1734) );
  OAI2B2X1 U6154 ( .A1N(Output1[10]), .A0(n2379), .B0(n4945), .B1(n2381), .Y(
        n1735) );
  CLKNAND2X2 U6155 ( .A(n3977), .B(n3734), .Y(n2381) );
  CLKINVX1 U6156 ( .A(dec), .Y(n3734) );
  CLKNAND2X2 U6157 ( .A(dec), .B(n3977), .Y(n2379) );
  XOR2X1 U6158 ( .A(n1952), .B(n4946), .Y(Output1[10]) );
  NOR2X1 U6159 ( .A(n254), .B(n4945), .Y(n4946) );
  CLKINVX1 U6160 ( .A(Input1[10]), .Y(n4945) );
  OAI221X1 U6161 ( .A0(n2136), .A1(n2274), .B0(n4881), .B1(n2273), .C0(n4947), 
        .Y(n1952) );
  MXI2X1 U6162 ( .A(n4948), .B(n4949), .S0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[8]), .Y(n4947) );
  OAI21X1 U6163 ( .A0(n4950), .A1(n280), .B0(n2267), .Y(n4949) );
  NOR2X1 U6164 ( .A(n2021), .B(n2140), .Y(n4950) );
  NOR3X1 U6165 ( .A(n274), .B(n2021), .C(n2140), .Y(n4948) );
  CLKINVX1 U6166 ( .A(n4590), .Y(n2140) );
  XNOR2X1 U6167 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_2_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[10]), .Y(n4590) );
  XOR2X1 U6168 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_3_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[11]), .Y(n2021) );
  XOR2X1 U6169 ( .A(n3918), .B(Inst_forkAE_CipherInst_RF_S_MID_C1[60]), .Y(
        n4881) );
  XNOR2X1 U6170 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[108]), .B(n4867), .Y(
        n3918) );
  XOR2X1 U6171 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[58]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_58_), .Y(n4867) );
  MXI2X1 U6172 ( .A(n4707), .B(n4951), .S0(n316), .Y(n2136) );
  XOR2X1 U6173 ( .A(Inst_forkAE_CipherInst_RF_S_MID_C1[20]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[116]), .Y(n4951) );
  XOR2X1 U6174 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_3_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_C1[12]), .Y(n4707) );
  OAI221X1 U6175 ( .A0(n1765), .A1(n165), .B0(n1968), .B1(n152), .C0(n4952), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_1_N3) );
  AOI22XL U6176 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_1_), 
        .B0(n219), .B1(Input1[1]), .Y(n4952) );
  AOI22XL U6177 ( .A0(Input1[1]), .A1(n2627), .B0(n1989), .B1(Output1[1]), .Y(
        n1765) );
  XOR2X1 U6178 ( .A(n4953), .B(n1968), .Y(Output1[1]) );
  CLKINVX1 U6179 ( .A(n4954), .Y(n1968) );
  OAI221X1 U6180 ( .A0(n2025), .A1(n2274), .B0(n3614), .B1(n2273), .C0(n4955), 
        .Y(n4954) );
  AOI22XL U6181 ( .A0(n291), .A1(n2049), .B0(
        Inst_forkAE_CipherInst_RF_S_MID_D1[3]), .B1(n300), .Y(n4955) );
  XOR2X1 U6182 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_1_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[3]), .Y(n2049) );
  XOR2X1 U6183 ( .A(n4041), .B(n4179), .Y(n3614) );
  CLKINVX1 U6184 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[55]), .Y(n4179) );
  XOR2X1 U6185 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[103]), .B(n4936), .Y(
        n4041) );
  XOR2X1 U6186 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[17]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_17_), .Y(n4936) );
  MXI2X1 U6187 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[7]), .B(n4956), .S0(
        n316), .Y(n2025) );
  XOR2X1 U6188 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[15]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[111]), .Y(n4956) );
  CLKNAND2X2 U6189 ( .A(Input1[1]), .B(n2288), .Y(n4953) );
  OAI221X1 U6190 ( .A0(n1768), .A1(n165), .B0(n1973), .B1(n152), .C0(n4957), 
        .Y(Inst_forkAE_CipherInst_RF_RS1_SFF_0_N3) );
  AOI22XL U6191 ( .A0(n190), .A1(Inst_forkAE_MainPart1_Tag_Reg_Output_0_), 
        .B0(n219), .B1(Input1[0]), .Y(n4957) );
  CLKINVX1 U6192 ( .A(n2302), .Y(n2249) );
  NOR2X1 U6193 ( .A(gen_tag), .B(a_data), .Y(n2000) );
  CLKINVX1 U6194 ( .A(n2300), .Y(n2248) );
  CLKNAND2X2 U6195 ( .A(n4958), .B(n145), .Y(n2300) );
  AOI22XL U6196 ( .A0(Input1[0]), .A1(n2627), .B0(n1989), .B1(Output1[0]), .Y(
        n1768) );
  XOR2X1 U6197 ( .A(n4959), .B(n1973), .Y(Output1[0]) );
  AOI221XL U6198 ( .A0(n3983), .A1(n297), .B0(n2166), .B1(n2293), .C0(n4960), 
        .Y(n1973) );
  AO22X1 U6199 ( .A0(n266), .A1(n3621), .B0(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]), .B1(n292), .Y(n4960) );
  CLKNAND2X2 U6200 ( .A(n2273), .B(n2244), .Y(n2266) );
  XOR2X1 U6201 ( .A(n2226), .B(n4051), .Y(n3621) );
  XNOR2X1 U6202 ( .A(n4933), .B(n3606), .Y(n4051) );
  XNOR2X1 U6203 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_24_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[98]), .Y(n3606) );
  XOR2X1 U6204 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[16]), .B(
        Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_16_), .Y(n4933) );
  CLKINVX1 U6205 ( .A(n4156), .Y(n2226) );
  XNOR2X1 U6206 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_12_), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[50]), .Y(n4156) );
  CLKINVX1 U6207 ( .A(n2273), .Y(n2260) );
  CLKINVX1 U6208 ( .A(n4226), .Y(n2166) );
  MXI2X1 U6209 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[1]), .B(n4961), .S0(
        n306), .Y(n4226) );
  XOR2X1 U6210 ( .A(Inst_forkAE_CipherInst_RF_S_MID_D1[9]), .B(
        Inst_forkAE_CipherInst_RF_S_MID_D1[105]), .Y(n4961) );
  CLKINVX1 U6211 ( .A(n2267), .Y(n2286) );
  XOR2X1 U6212 ( .A(Inst_forkAE_CipherInst_RF_STATE_EX1_0_), .B(
        Inst_forkAE_CipherInst_RF_SHIFT1_OUT[15]), .Y(n3983) );
  CLKNAND2X2 U6213 ( .A(Input1[0]), .B(n2288), .Y(n4959) );
  NOR2X1 U6214 ( .A(n2288), .B(dec), .Y(n2627) );
  OAI221X1 U6215 ( .A0(n335), .A1(n4962), .B0(n355), .B1(n4964), .C0(n4965), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_99_N3) );
  OAI221X1 U6216 ( .A0(n332), .A1(n4966), .B0(n364), .B1(n4967), .C0(n4968), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_98_N3) );
  OAI221X1 U6217 ( .A0(n332), .A1(n4969), .B0(n364), .B1(n4970), .C0(n4971), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_97_N3) );
  OAI221X1 U6218 ( .A0(n4972), .A1(n336), .B0(n364), .B1(n4973), .C0(n4974), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_96_N3) );
  XOR2X1 U6219 ( .A(n4975), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_87_), 
        .Y(n4972) );
  OAI221X1 U6220 ( .A0(n332), .A1(n4976), .B0(n364), .B1(n4977), .C0(n4978), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_95_N3) );
  CLKINVX1 U6221 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_95_), .Y(n4977) );
  OAI221X1 U6222 ( .A0(n332), .A1(n4979), .B0(n364), .B1(n4980), .C0(n4981), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_94_N3) );
  OAI221X1 U6223 ( .A0(n332), .A1(n4982), .B0(n364), .B1(n4983), .C0(n4984), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_93_N3) );
  OAI221X1 U6224 ( .A0(n332), .A1(n4985), .B0(n364), .B1(n4986), .C0(n4987), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_92_N3) );
  OAI221X1 U6225 ( .A0(n333), .A1(n4988), .B0(n364), .B1(n4989), .C0(n4990), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_91_N3) );
  OAI221X1 U6226 ( .A0(n332), .A1(n4991), .B0(n363), .B1(n4992), .C0(n4993), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_90_N3) );
  OAI221X1 U6227 ( .A0(n3054), .A1(n336), .B0(n2956), .B1(n370), .C0(n4994), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_9_N3) );
  OAI221X1 U6228 ( .A0(n335), .A1(n4995), .B0(n364), .B1(n4996), .C0(n4997), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_89_N3) );
  OAI221X1 U6229 ( .A0(n4998), .A1(n337), .B0(n363), .B1(n4999), .C0(n5000), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_88_N3) );
  XOR2X1 U6230 ( .A(n4979), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_111_), 
        .Y(n4998) );
  OAI221X1 U6231 ( .A0(n335), .A1(n5001), .B0(n364), .B1(n5002), .C0(n5003), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_87_N3) );
  CLKINVX1 U6232 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_87_), .Y(n5002) );
  OAI221X1 U6233 ( .A0(n334), .A1(n5004), .B0(n362), .B1(n5005), .C0(n5006), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_86_N3) );
  OAI221X1 U6234 ( .A0(n335), .A1(n5007), .B0(n364), .B1(n4975), .C0(n5008), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_85_N3) );
  OAI221X1 U6235 ( .A0(n335), .A1(n5009), .B0(n363), .B1(n5010), .C0(n5011), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_84_N3) );
  OAI221X1 U6236 ( .A0(n334), .A1(n5012), .B0(n364), .B1(n5013), .C0(n5014), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_83_N3) );
  OAI221X1 U6237 ( .A0(n334), .A1(n5015), .B0(n4962), .B1(n370), .C0(n5016), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_82_N3) );
  CLKINVX1 U6238 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_82_), .Y(n4962) );
  OAI221X1 U6239 ( .A0(n335), .A1(n5017), .B0(n363), .B1(n4966), .C0(n5018), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_81_N3) );
  CLKINVX1 U6240 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_81_), .Y(n4966) );
  OAI221X1 U6241 ( .A0(n5019), .A1(n337), .B0(n363), .B1(n4969), .C0(n5020), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_80_N3) );
  CLKINVX1 U6242 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_80_), .Y(n4969) );
  XOR2X1 U6243 ( .A(n5004), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_79_), 
        .Y(n5019) );
  OAI221X1 U6244 ( .A0(n2543), .A1(n337), .B0(n2964), .B1(n371), .C0(n5021), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_8_N3) );
  OAI221X1 U6245 ( .A0(n334), .A1(n4980), .B0(n363), .B1(n5022), .C0(n5023), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_79_N3) );
  CLKINVX1 U6246 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_79_), .Y(n5022) );
  CLKINVX1 U6247 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_94_), .Y(n4980) );
  OAI221X1 U6248 ( .A0(n334), .A1(n4983), .B0(n363), .B1(n5001), .C0(n5024), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_78_N3) );
  CLKINVX1 U6249 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_78_), .Y(n5001) );
  OAI221X1 U6250 ( .A0(n335), .A1(n4986), .B0(n363), .B1(n5004), .C0(n5025), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_77_N3) );
  CLKINVX1 U6251 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_77_), .Y(n5004) );
  CLKINVX1 U6252 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_92_), .Y(n4986) );
  OAI221X1 U6253 ( .A0(n334), .A1(n4989), .B0(n363), .B1(n5007), .C0(n5026), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_76_N3) );
  CLKINVX1 U6254 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_76_), .Y(n5007) );
  CLKINVX1 U6255 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_91_), .Y(n4989) );
  OAI221X1 U6256 ( .A0(n333), .A1(n4992), .B0(n362), .B1(n5009), .C0(n5027), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_75_N3) );
  CLKINVX1 U6257 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_75_), .Y(n5009) );
  CLKINVX1 U6258 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_90_), .Y(n4992) );
  OAI221X1 U6259 ( .A0(n334), .A1(n4996), .B0(n363), .B1(n5012), .C0(n5028), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_74_N3) );
  CLKINVX1 U6260 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_74_), .Y(n5012) );
  CLKINVX1 U6261 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_89_), .Y(n4996) );
  OAI221X1 U6262 ( .A0(n334), .A1(n4999), .B0(n362), .B1(n5015), .C0(n5029), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_73_N3) );
  CLKINVX1 U6263 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_73_), .Y(n5015) );
  CLKINVX1 U6264 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_88_), .Y(n4999) );
  OAI221X1 U6265 ( .A0(n5030), .A1(n337), .B0(n363), .B1(n5017), .C0(n5031), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_72_N3) );
  CLKINVX1 U6266 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_72_), .Y(n5017) );
  XOR2X1 U6267 ( .A(n4983), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_95_), 
        .Y(n5030) );
  CLKINVX1 U6268 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_93_), .Y(n4983) );
  OAI221X1 U6269 ( .A0(n332), .A1(n5032), .B0(n362), .B1(n5033), .C0(n5034), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_71_N3) );
  CLKINVX1 U6270 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_71_), .Y(n5033) );
  OAI221X1 U6271 ( .A0(n332), .A1(n5035), .B0(n363), .B1(n5036), .C0(n5037), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_70_N3) );
  OAI221X1 U6272 ( .A0(n5038), .A1(n365), .B0(n5039), .B1(n337), .C0(n5040), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_7_N3) );
  XOR2X1 U6273 ( .A(n3382), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_6_), 
        .Y(n5038) );
  OAI221X1 U6274 ( .A0(n332), .A1(n5041), .B0(n363), .B1(n5042), .C0(n5043), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_69_N3) );
  OAI221X1 U6275 ( .A0(n332), .A1(n4964), .B0(n362), .B1(n5044), .C0(n5045), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_68_N3) );
  CLKINVX1 U6276 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_99_), .Y(n4964) );
  OAI221X1 U6277 ( .A0(n331), .A1(n4967), .B0(n362), .B1(n5046), .C0(n5047), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_67_N3) );
  CLKINVX1 U6278 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_98_), .Y(n4967) );
  OAI221X1 U6279 ( .A0(n331), .A1(n4970), .B0(n362), .B1(n5048), .C0(n5049), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_66_N3) );
  CLKINVX1 U6280 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_97_), .Y(n4970) );
  OAI221X1 U6281 ( .A0(n331), .A1(n4973), .B0(n362), .B1(n5050), .C0(n5051), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_65_N3) );
  CLKINVX1 U6282 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_96_), .Y(n4973) );
  OAI221X1 U6283 ( .A0(n5052), .A1(n336), .B0(n362), .B1(n5053), .C0(n5054), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_64_N3) );
  XOR2X1 U6284 ( .A(n5035), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_103_), 
        .Y(n5052) );
  OAI221X1 U6285 ( .A0(n5055), .A1(n365), .B0(n3276), .B1(n338), .C0(n5056), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_63_N3) );
  XOR2X1 U6286 ( .A(n3474), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_62_), 
        .Y(n5055) );
  OAI221X1 U6287 ( .A0(n3288), .A1(n340), .B0(n3440), .B1(n372), .C0(n5057), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_62_N3) );
  OAI221X1 U6288 ( .A0(n3294), .A1(n340), .B0(n3452), .B1(n372), .C0(n5058), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_61_N3) );
  OAI221X1 U6289 ( .A0(n3287), .A1(n340), .B0(n3470), .B1(n372), .C0(n5059), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_60_N3) );
  OAI221X1 U6290 ( .A0(n5060), .A1(n340), .B0(n3358), .B1(n372), .C0(n5061), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_6_N3) );
  OAI221X1 U6291 ( .A0(n3314), .A1(n340), .B0(n3451), .B1(n372), .C0(n5062), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_59_N3) );
  OAI221X1 U6292 ( .A0(n3327), .A1(n339), .B0(n3492), .B1(n372), .C0(n5063), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_58_N3) );
  OAI221X1 U6293 ( .A0(n5064), .A1(n339), .B0(n3572), .B1(n372), .C0(n5065), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_57_N3) );
  OAI221X1 U6294 ( .A0(n3298), .A1(n339), .B0(n5066), .B1(n372), .C0(n5067), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_56_N3) );
  OAI221X1 U6295 ( .A0(n5068), .A1(n365), .B0(n3358), .B1(n345), .C0(n5069), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_55_N3) );
  CLKINVX1 U6296 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_7_), .Y(n3358)
         );
  XOR2X1 U6297 ( .A(n3298), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_54_), 
        .Y(n5068) );
  CLKINVX1 U6298 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_48_), .Y(n3298) );
  OAI221X1 U6299 ( .A0(n3371), .A1(n339), .B0(n3276), .B1(n372), .C0(n5070), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_54_N3) );
  CLKINVX1 U6300 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_55_), .Y(n3276) );
  OAI221X1 U6301 ( .A0(n3378), .A1(n339), .B0(n3288), .B1(n373), .C0(n5071), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_53_N3) );
  CLKINVX1 U6302 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_54_), .Y(n3288) );
  OAI221X1 U6303 ( .A0(n3370), .A1(n339), .B0(n3294), .B1(n373), .C0(n5072), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_52_N3) );
  CLKINVX1 U6304 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_53_), .Y(n3294) );
  OAI221X1 U6305 ( .A0(n3400), .A1(n339), .B0(n3287), .B1(n373), .C0(n5073), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_51_N3) );
  CLKINVX1 U6306 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_52_), .Y(n3287) );
  OAI221X1 U6307 ( .A0(n3414), .A1(n339), .B0(n3314), .B1(n373), .C0(n5074), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_50_N3) );
  CLKINVX1 U6308 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_51_), .Y(n3314) );
  OAI221X1 U6309 ( .A0(n2736), .A1(n339), .B0(n3371), .B1(n373), .C0(n5075), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_5_N3) );
  CLKINVX1 U6310 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_6_), .Y(n3371)
         );
  OAI221X1 U6311 ( .A0(n5076), .A1(n339), .B0(n3327), .B1(n373), .C0(n5077), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_49_N3) );
  CLKINVX1 U6312 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_50_), .Y(n3327) );
  OAI221X1 U6313 ( .A0(n3382), .A1(n339), .B0(n5064), .B1(n373), .C0(n5078), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_48_N3) );
  CLKINVX1 U6314 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_49_), .Y(n5064) );
  CLKINVX1 U6315 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_0_), .Y(n3382)
         );
  OAI221X1 U6316 ( .A0(n5079), .A1(n365), .B0(n3440), .B1(n345), .C0(n5080), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_47_N3) );
  CLKINVX1 U6317 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_63_), .Y(n3440) );
  XOR2X1 U6318 ( .A(n2341), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_), 
        .Y(n5079) );
  OAI221X1 U6319 ( .A0(n3452), .A1(n339), .B0(n5081), .B1(n373), .C0(n5082), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_46_N3) );
  CLKINVX1 U6320 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_62_), .Y(n3452) );
  OAI221X1 U6321 ( .A0(n3470), .A1(n339), .B0(n5083), .B1(n373), .C0(n5084), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_45_N3) );
  CLKINVX1 U6322 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_61_), .Y(n3470) );
  OAI221X1 U6323 ( .A0(n3451), .A1(n338), .B0(n2830), .B1(n373), .C0(n5085), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_44_N3) );
  CLKINVX1 U6324 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_60_), .Y(n3451) );
  OAI221X1 U6325 ( .A0(n3492), .A1(n338), .B0(n2328), .B1(n373), .C0(n5086), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_43_N3) );
  CLKINVX1 U6326 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_59_), .Y(n3492) );
  OAI221X1 U6327 ( .A0(n3572), .A1(n338), .B0(n5087), .B1(n373), .C0(n5088), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_42_N3) );
  CLKINVX1 U6328 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_58_), .Y(n3572) );
  OAI221X1 U6329 ( .A0(n5066), .A1(n338), .B0(n2861), .B1(n374), .C0(n5089), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_41_N3) );
  CLKINVX1 U6330 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_57_), .Y(n5066) );
  OAI221X1 U6331 ( .A0(n3474), .A1(n338), .B0(n2880), .B1(n374), .C0(n5090), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_40_N3) );
  CLKINVX1 U6332 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_56_), .Y(n3474) );
  OAI221X1 U6333 ( .A0(n2623), .A1(n338), .B0(n3378), .B1(n374), .C0(n5091), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_4_N3) );
  CLKINVX1 U6334 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_5_), .Y(n3378)
         );
  OAI221X1 U6335 ( .A0(n5092), .A1(n365), .B0(n5093), .B1(n343), .C0(n5094), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_39_N3) );
  XOR2X1 U6336 ( .A(n2646), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_), 
        .Y(n5092) );
  OAI221X1 U6337 ( .A0(n3543), .A1(n338), .B0(n5039), .B1(n374), .C0(n5095), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_38_N3) );
  CLKINVX1 U6338 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_39_), .Y(n5039) );
  OAI221X1 U6339 ( .A0(n3550), .A1(n338), .B0(n5060), .B1(n374), .C0(n5096), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_37_N3) );
  CLKINVX1 U6340 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_38_), .Y(n5060) );
  OAI221X1 U6341 ( .A0(n3539), .A1(n338), .B0(n2736), .B1(n374), .C0(n5097), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_36_N3) );
  CLKINVX1 U6342 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_37_), .Y(n2736) );
  OAI221X1 U6343 ( .A0(n5098), .A1(n338), .B0(n2623), .B1(n374), .C0(n5099), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_35_N3) );
  CLKINVX1 U6344 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_36_), .Y(n2623) );
  OAI221X1 U6345 ( .A0(n3198), .A1(n338), .B0(n5100), .B1(n374), .C0(n5101), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_34_N3) );
  OAI221X1 U6346 ( .A0(n5102), .A1(n338), .B0(n2778), .B1(n374), .C0(n5103), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_33_N3) );
  OAI221X1 U6347 ( .A0(n3555), .A1(n338), .B0(n2787), .B1(n374), .C0(n5104), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_32_N3) );
  OAI221X1 U6348 ( .A0(n5105), .A1(n365), .B0(n5081), .B1(n345), .C0(n5106), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_31_N3) );
  CLKINVX1 U6349 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_47_), .Y(n5081) );
  XOR2X1 U6350 ( .A(n2543), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_), 
        .Y(n5105) );
  CLKINVX1 U6351 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_24_), .Y(n2543) );
  OAI221X1 U6352 ( .A0(n5083), .A1(n337), .B0(n5107), .B1(n374), .C0(n5108), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_30_N3) );
  CLKINVX1 U6353 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_46_), .Y(n5083) );
  OAI221X1 U6354 ( .A0(n5100), .A1(n337), .B0(n3370), .B1(n374), .C0(n5109), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_3_N3) );
  CLKINVX1 U6355 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_4_), .Y(n3370)
         );
  CLKINVX1 U6356 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_35_), .Y(n5100) );
  OAI221X1 U6357 ( .A0(n2830), .A1(n337), .B0(n5110), .B1(n375), .C0(n5111), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_29_N3) );
  CLKINVX1 U6358 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_45_), .Y(n2830) );
  OAI221X1 U6359 ( .A0(n2328), .A1(n337), .B0(n3016), .B1(n375), .C0(n5112), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_28_N3) );
  CLKINVX1 U6360 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_44_), .Y(n2328) );
  OAI221X1 U6361 ( .A0(n5087), .A1(n337), .B0(n2531), .B1(n375), .C0(n5113), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_27_N3) );
  CLKINVX1 U6362 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_43_), .Y(n5087) );
  OAI221X1 U6363 ( .A0(n2861), .A1(n337), .B0(n5114), .B1(n375), .C0(n5115), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_26_N3) );
  CLKINVX1 U6364 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_42_), .Y(n2861) );
  OAI221X1 U6365 ( .A0(n2880), .A1(n336), .B0(n3046), .B1(n375), .C0(n5116), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_25_N3) );
  CLKINVX1 U6366 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_41_), .Y(n2880) );
  OAI221X1 U6367 ( .A0(n2341), .A1(n336), .B0(n3054), .B1(n375), .C0(n5117), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_24_N3) );
  CLKINVX1 U6368 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_25_), .Y(n3054) );
  CLKINVX1 U6369 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_40_), .Y(n2341) );
  OAI221X1 U6370 ( .A0(n5118), .A1(n365), .B0(n5119), .B1(n345), .C0(n5120), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_23_N3) );
  XOR2X1 U6371 ( .A(n3555), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_22_), 
        .Y(n5118) );
  CLKINVX1 U6372 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_16_), .Y(n3555) );
  OAI221X1 U6373 ( .A0(n5121), .A1(n337), .B0(n5093), .B1(n375), .C0(n5122), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_22_N3) );
  CLKINVX1 U6374 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_23_), .Y(n5093) );
  OAI221X1 U6375 ( .A0(n2926), .A1(n336), .B0(n3543), .B1(n375), .C0(n5123), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_21_N3) );
  CLKINVX1 U6376 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_22_), .Y(n3543) );
  OAI221X1 U6377 ( .A0(n2430), .A1(n336), .B0(n3550), .B1(n375), .C0(n5124), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_20_N3) );
  CLKINVX1 U6378 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_21_), .Y(n3550) );
  OAI221X1 U6379 ( .A0(n2778), .A1(n336), .B0(n3400), .B1(n375), .C0(n5125), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_2_N3) );
  CLKINVX1 U6380 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_3_), .Y(n3400)
         );
  CLKINVX1 U6381 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_34_), .Y(n2778) );
  OAI221X1 U6382 ( .A0(n5126), .A1(n336), .B0(n3539), .B1(n375), .C0(n5127), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_19_N3) );
  CLKINVX1 U6383 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_20_), .Y(n3539) );
  OAI221X1 U6384 ( .A0(n2956), .A1(n336), .B0(n5098), .B1(n375), .C0(n5128), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_18_N3) );
  CLKINVX1 U6385 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_19_), .Y(n5098) );
  CLKINVX1 U6386 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_10_), .Y(n2956) );
  OAI221X1 U6387 ( .A0(n2964), .A1(n336), .B0(n3198), .B1(n375), .C0(n5129), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_17_N3) );
  CLKINVX1 U6388 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_18_), .Y(n3198) );
  CLKINVX1 U6389 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_9_), .Y(n2964)
         );
  OAI221X1 U6390 ( .A0(n2442), .A1(n337), .B0(n5102), .B1(n375), .C0(n5130), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_16_N3) );
  CLKINVX1 U6391 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_17_), .Y(n5102) );
  CLKINVX1 U6392 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_8_), .Y(n2442)
         );
  OAI221X1 U6393 ( .A0(n5131), .A1(n365), .B0(n5107), .B1(n345), .C0(n5132), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_15_N3) );
  CLKINVX1 U6394 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_31_), .Y(n5107) );
  XOR2X1 U6395 ( .A(n5121), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_8_), 
        .Y(n5131) );
  OAI221X1 U6396 ( .A0(n5110), .A1(n340), .B0(n5119), .B1(n376), .C0(n5133), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_14_N3) );
  CLKINVX1 U6397 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_15_), .Y(n5119) );
  CLKINVX1 U6398 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_30_), .Y(n5110) );
  OAI221X1 U6399 ( .A0(n3016), .A1(n340), .B0(n5121), .B1(n376), .C0(n5134), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_13_N3) );
  CLKINVX1 U6400 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_14_), .Y(n5121) );
  CLKINVX1 U6401 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_29_), .Y(n3016) );
  OAI221X1 U6402 ( .A0(n327), .A1(n5135), .B0(n362), .B1(n5136), .C0(n5137), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_127_N3) );
  CLKINVX1 U6403 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_127_), .Y(
        n5136) );
  OAI221X1 U6404 ( .A0(n327), .A1(n5138), .B0(n362), .B1(n5139), .C0(n5140), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_126_N3) );
  OAI221X1 U6405 ( .A0(n327), .A1(n5141), .B0(n362), .B1(n5142), .C0(n5143), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_125_N3) );
  OAI221X1 U6406 ( .A0(n327), .A1(n5144), .B0(n362), .B1(n5145), .C0(n5146), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_124_N3) );
  OAI221X1 U6407 ( .A0(n327), .A1(n5147), .B0(n361), .B1(n5148), .C0(n5149), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_123_N3) );
  OAI221X1 U6408 ( .A0(n327), .A1(n5150), .B0(n360), .B1(n5151), .C0(n5152), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_122_N3) );
  OAI221X1 U6409 ( .A0(n328), .A1(n5153), .B0(n359), .B1(n5154), .C0(n5155), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_121_N3) );
  OAI221X1 U6410 ( .A0(n5156), .A1(n340), .B0(n359), .B1(n5157), .C0(n5158), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_120_N3) );
  XOR2X1 U6411 ( .A(n5138), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_119_), 
        .Y(n5156) );
  OAI221X1 U6412 ( .A0(n2531), .A1(n340), .B0(n2926), .B1(n376), .C0(n5159), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_12_N3) );
  CLKINVX1 U6413 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_13_), .Y(n2926) );
  CLKINVX1 U6414 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_28_), .Y(n2531) );
  OAI221X1 U6415 ( .A0(n328), .A1(n5036), .B0(n359), .B1(n5160), .C0(n5161), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_119_N3) );
  CLKINVX1 U6416 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_119_), .Y(
        n5160) );
  CLKINVX1 U6417 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_70_), .Y(n5036) );
  OAI221X1 U6418 ( .A0(n328), .A1(n5042), .B0(n359), .B1(n5135), .C0(n5162), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_118_N3) );
  CLKINVX1 U6419 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_118_), .Y(
        n5135) );
  OAI221X1 U6420 ( .A0(n328), .A1(n5044), .B0(n359), .B1(n5138), .C0(n5163), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_117_N3) );
  CLKINVX1 U6421 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_117_), .Y(
        n5138) );
  CLKINVX1 U6422 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_68_), .Y(n5044) );
  OAI221X1 U6423 ( .A0(n328), .A1(n5046), .B0(n359), .B1(n5141), .C0(n5164), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_116_N3) );
  CLKINVX1 U6424 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_116_), .Y(
        n5141) );
  CLKINVX1 U6425 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_67_), .Y(n5046) );
  OAI221X1 U6426 ( .A0(n328), .A1(n5048), .B0(n359), .B1(n5144), .C0(n5165), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_115_N3) );
  CLKINVX1 U6427 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_115_), .Y(
        n5144) );
  CLKINVX1 U6428 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_66_), .Y(n5048) );
  OAI221X1 U6429 ( .A0(n328), .A1(n5050), .B0(n359), .B1(n5147), .C0(n5166), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_114_N3) );
  CLKINVX1 U6430 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_114_), .Y(
        n5147) );
  CLKINVX1 U6431 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_65_), .Y(n5050) );
  OAI221X1 U6432 ( .A0(n328), .A1(n5053), .B0(n358), .B1(n5150), .C0(n5167), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_113_N3) );
  CLKINVX1 U6433 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_113_), .Y(
        n5150) );
  CLKINVX1 U6434 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_64_), .Y(n5053) );
  OAI221X1 U6435 ( .A0(n5168), .A1(n340), .B0(n358), .B1(n5153), .C0(n5169), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_112_N3) );
  CLKINVX1 U6436 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_112_), .Y(
        n5153) );
  XOR2X1 U6437 ( .A(n5042), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_71_), 
        .Y(n5168) );
  CLKINVX1 U6438 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_69_), .Y(n5042) );
  OAI221X1 U6439 ( .A0(n328), .A1(n5139), .B0(n358), .B1(n5170), .C0(n5171), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_111_N3) );
  CLKINVX1 U6440 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_111_), .Y(
        n5170) );
  CLKINVX1 U6441 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_126_), .Y(
        n5139) );
  OAI221X1 U6442 ( .A0(n328), .A1(n5142), .B0(n358), .B1(n4976), .C0(n5172), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_110_N3) );
  CLKINVX1 U6443 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_110_), .Y(
        n4976) );
  OAI221X1 U6444 ( .A0(n5114), .A1(n340), .B0(n2430), .B1(n377), .C0(n5173), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_11_N3) );
  CLKINVX1 U6445 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_12_), .Y(n2430) );
  CLKINVX1 U6446 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_27_), .Y(n5114) );
  OAI221X1 U6447 ( .A0(n328), .A1(n5145), .B0(n358), .B1(n4979), .C0(n5174), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_109_N3) );
  CLKINVX1 U6448 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_109_), .Y(
        n4979) );
  CLKINVX1 U6449 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_124_), .Y(
        n5145) );
  OAI221X1 U6450 ( .A0(n328), .A1(n5148), .B0(n358), .B1(n4982), .C0(n5175), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_108_N3) );
  CLKINVX1 U6451 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_108_), .Y(
        n4982) );
  CLKINVX1 U6452 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_123_), .Y(
        n5148) );
  OAI221X1 U6453 ( .A0(n328), .A1(n5151), .B0(n358), .B1(n4985), .C0(n5176), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_107_N3) );
  CLKINVX1 U6454 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_107_), .Y(
        n4985) );
  CLKINVX1 U6455 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_122_), .Y(
        n5151) );
  OAI221X1 U6456 ( .A0(n329), .A1(n5154), .B0(n358), .B1(n4988), .C0(n5177), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_106_N3) );
  CLKINVX1 U6457 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_106_), .Y(
        n4988) );
  CLKINVX1 U6458 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_121_), .Y(
        n5154) );
  OAI221X1 U6459 ( .A0(n329), .A1(n5157), .B0(n358), .B1(n4991), .C0(n5178), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_105_N3) );
  CLKINVX1 U6460 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_105_), .Y(
        n4991) );
  CLKINVX1 U6461 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_120_), .Y(
        n5157) );
  OAI221X1 U6462 ( .A0(n5179), .A1(n340), .B0(n358), .B1(n4995), .C0(n5180), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_104_N3) );
  CLKINVX1 U6463 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_104_), .Y(
        n4995) );
  XOR2X1 U6464 ( .A(n5142), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_127_), 
        .Y(n5179) );
  CLKINVX1 U6465 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_125_), .Y(
        n5142) );
  OAI221X1 U6466 ( .A0(n329), .A1(n5005), .B0(n358), .B1(n5181), .C0(n5182), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_103_N3) );
  CLKINVX1 U6467 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_103_), .Y(
        n5181) );
  CLKINVX1 U6468 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_86_), .Y(n5005) );
  OAI221X1 U6469 ( .A0(n329), .A1(n4975), .B0(n358), .B1(n5032), .C0(n5183), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_102_N3) );
  CLKINVX1 U6470 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_102_), .Y(
        n5032) );
  CLKINVX1 U6471 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_85_), .Y(n4975) );
  OAI221X1 U6472 ( .A0(n329), .A1(n5010), .B0(n358), .B1(n5035), .C0(n5184), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_101_N3) );
  CLKINVX1 U6473 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_101_), .Y(
        n5035) );
  CLKINVX1 U6474 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_84_), .Y(n5010) );
  OAI221X1 U6475 ( .A0(n329), .A1(n5013), .B0(n357), .B1(n5041), .C0(n5185), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_100_N3) );
  CLKINVX1 U6476 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_100_), .Y(
        n5041) );
  CLKINVX1 U6477 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_83_), .Y(n5013) );
  OAI221X1 U6478 ( .A0(n3046), .A1(n341), .B0(n5126), .B1(n373), .C0(n5186), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_10_N3) );
  CLKINVX1 U6479 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_11_), .Y(n5126) );
  CLKINVX1 U6480 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_26_), .Y(n3046) );
  OAI221X1 U6481 ( .A0(n2787), .A1(n341), .B0(n3414), .B1(n372), .C0(n5187), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_1_N3) );
  CLKINVX1 U6482 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_2_), .Y(n3414)
         );
  CLKINVX1 U6483 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_33_), .Y(n2787) );
  OAI221X1 U6484 ( .A0(n2646), .A1(n341), .B0(n5076), .B1(n372), .C0(n5188), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_2_SFF_0_N3) );
  CLKINVX1 U6485 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_1_), .Y(n5076)
         );
  CLKINVX1 U6486 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_2_Inv_32_), .Y(n2646) );
  OAI221X1 U6487 ( .A0(n329), .A1(n5189), .B0(n357), .B1(n5190), .C0(n4965), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_99_N3) );
  AOI22XL U6488 ( .A0(n5191), .A1(n414), .B0(n398), .B1(K1[99]), .Y(n4965) );
  OAI221X1 U6489 ( .A0(n329), .A1(n5193), .B0(n357), .B1(n5194), .C0(n4968), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_98_N3) );
  AOI22XL U6490 ( .A0(n5195), .A1(n414), .B0(n396), .B1(K1[98]), .Y(n4968) );
  OAI221X1 U6491 ( .A0(n329), .A1(n5196), .B0(n357), .B1(n5197), .C0(n4971), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_97_N3) );
  AOI22XL U6492 ( .A0(K1[39]), .A1(n414), .B0(n396), .B1(K1[97]), .Y(n4971) );
  OAI221X1 U6493 ( .A0(n5198), .A1(n341), .B0(n357), .B1(n5199), .C0(n4974), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_96_N3) );
  AOI22XL U6494 ( .A0(n414), .A1(K1[38]), .B0(n396), .B1(K1[96]), .Y(n4974) );
  XOR2X1 U6495 ( .A(n5200), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_87_), 
        .Y(n5198) );
  OAI221X1 U6496 ( .A0(n329), .A1(n5201), .B0(n357), .B1(n5202), .C0(n4978), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_95_N3) );
  AOI2BB2X1 U6497 ( .B0(n389), .B1(K1[95]), .A0N(n5203), .A1N(n409), .Y(n4978)
         );
  XOR2X1 U6498 ( .A(n5204), .B(K1[29]), .Y(n5203) );
  CLKINVX1 U6499 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_95_), .Y(n5202) );
  OAI221X1 U6500 ( .A0(n329), .A1(n5205), .B0(n357), .B1(n5206), .C0(n4981), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_94_N3) );
  AOI2BB2X1 U6501 ( .B0(n389), .B1(K1[94]), .A0N(n5207), .A1N(n409), .Y(n4981)
         );
  XOR2X1 U6502 ( .A(n5208), .B(K1[28]), .Y(n5207) );
  OAI221X1 U6503 ( .A0(n329), .A1(n5209), .B0(n357), .B1(n5210), .C0(n4984), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_93_N3) );
  AOI2BB2X1 U6504 ( .B0(n389), .B1(K1[93]), .A0N(n5204), .A1N(n410), .Y(n4984)
         );
  XNOR2X1 U6505 ( .A(K1[27]), .B(n5211), .Y(n5204) );
  OAI221X1 U6506 ( .A0(n329), .A1(n5212), .B0(n357), .B1(n5213), .C0(n4987), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_92_N3) );
  AOI2BB2X1 U6507 ( .B0(n389), .B1(K1[92]), .A0N(n5208), .A1N(n408), .Y(n4987)
         );
  XNOR2X1 U6508 ( .A(K1[26]), .B(n5214), .Y(n5208) );
  OAI221X1 U6509 ( .A0(n330), .A1(n5215), .B0(n357), .B1(n5216), .C0(n4990), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_91_N3) );
  AOI22XL U6510 ( .A0(n5211), .A1(n414), .B0(n397), .B1(K1[91]), .Y(n4990) );
  XOR2X1 U6511 ( .A(K1[31]), .B(K1[25]), .Y(n5211) );
  OAI221X1 U6512 ( .A0(n330), .A1(n5217), .B0(n357), .B1(n5218), .C0(n4993), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_90_N3) );
  AOI22XL U6513 ( .A0(n5214), .A1(n414), .B0(n397), .B1(K1[90]), .Y(n4993) );
  XOR2X1 U6514 ( .A(K1[30]), .B(K1[24]), .Y(n5214) );
  OAI221X1 U6515 ( .A0(n5219), .A1(n341), .B0(n5220), .B1(n371), .C0(n4994), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_9_N3) );
  AOI2BB2X1 U6516 ( .B0(n389), .B1(K1[9]), .A0N(n5221), .A1N(n409), .Y(n4994)
         );
  XOR2X1 U6517 ( .A(K1[80]), .B(n5222), .Y(n5221) );
  OAI221X1 U6518 ( .A0(n330), .A1(n5223), .B0(n357), .B1(n5224), .C0(n4997), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_89_N3) );
  AOI22XL U6519 ( .A0(n414), .A1(K1[31]), .B0(n397), .B1(K1[89]), .Y(n4997) );
  OAI221X1 U6520 ( .A0(n5225), .A1(n341), .B0(n357), .B1(n5226), .C0(n5000), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_88_N3) );
  AOI22XL U6521 ( .A0(n414), .A1(K1[30]), .B0(n397), .B1(K1[88]), .Y(n5000) );
  XOR2X1 U6522 ( .A(n5205), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_111_), 
        .Y(n5225) );
  OAI221X1 U6523 ( .A0(n330), .A1(n5227), .B0(n356), .B1(n5228), .C0(n5003), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_87_N3) );
  AOI2BB2X1 U6524 ( .B0(n389), .B1(K1[87]), .A0N(n5229), .A1N(n410), .Y(n5003)
         );
  XOR2X1 U6525 ( .A(n5230), .B(K1[21]), .Y(n5229) );
  CLKINVX1 U6526 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_87_), .Y(n5228) );
  OAI221X1 U6527 ( .A0(n330), .A1(n5231), .B0(n356), .B1(n5232), .C0(n5006), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_86_N3) );
  AOI2BB2X1 U6528 ( .B0(n389), .B1(K1[86]), .A0N(n5233), .A1N(n408), .Y(n5006)
         );
  XOR2X1 U6529 ( .A(n5234), .B(K1[20]), .Y(n5233) );
  OAI221X1 U6530 ( .A0(n330), .A1(n5235), .B0(n356), .B1(n5200), .C0(n5008), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_85_N3) );
  AOI2BB2X1 U6531 ( .B0(n389), .B1(K1[85]), .A0N(n5230), .A1N(n409), .Y(n5008)
         );
  XNOR2X1 U6532 ( .A(K1[19]), .B(n5236), .Y(n5230) );
  OAI221X1 U6533 ( .A0(n332), .A1(n5237), .B0(n356), .B1(n5238), .C0(n5011), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_84_N3) );
  AOI2BB2X1 U6534 ( .B0(n389), .B1(K1[84]), .A0N(n5234), .A1N(n410), .Y(n5011)
         );
  XNOR2X1 U6535 ( .A(K1[18]), .B(n5239), .Y(n5234) );
  OAI221X1 U6536 ( .A0(n330), .A1(n5240), .B0(n356), .B1(n5241), .C0(n5014), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_83_N3) );
  AOI22XL U6537 ( .A0(n5236), .A1(n414), .B0(n397), .B1(K1[83]), .Y(n5014) );
  XOR2X1 U6538 ( .A(K1[23]), .B(K1[17]), .Y(n5236) );
  OAI221X1 U6539 ( .A0(n330), .A1(n5242), .B0(n356), .B1(n5189), .C0(n5016), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_82_N3) );
  AOI22XL U6540 ( .A0(n5239), .A1(n414), .B0(n397), .B1(K1[82]), .Y(n5016) );
  XOR2X1 U6541 ( .A(K1[22]), .B(K1[16]), .Y(n5239) );
  CLKINVX1 U6542 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_82_), .Y(n5189) );
  OAI221X1 U6543 ( .A0(n330), .A1(n5243), .B0(n356), .B1(n5193), .C0(n5018), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_81_N3) );
  AOI22XL U6544 ( .A0(n414), .A1(K1[23]), .B0(n398), .B1(K1[81]), .Y(n5018) );
  CLKINVX1 U6545 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_81_), .Y(n5193) );
  OAI221X1 U6546 ( .A0(n5244), .A1(n341), .B0(n356), .B1(n5196), .C0(n5020), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_80_N3) );
  AOI22XL U6547 ( .A0(n414), .A1(K1[22]), .B0(n397), .B1(K1[80]), .Y(n5020) );
  CLKINVX1 U6548 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_80_), .Y(n5196) );
  XOR2X1 U6549 ( .A(n5231), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_79_), 
        .Y(n5244) );
  OAI221X1 U6550 ( .A0(n5245), .A1(n341), .B0(n5246), .B1(n370), .C0(n5021), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_8_N3) );
  AOI22XL U6551 ( .A0(n414), .A1(K1[87]), .B0(n398), .B1(K1[8]), .Y(n5021) );
  OAI221X1 U6552 ( .A0(n330), .A1(n5206), .B0(n356), .B1(n5247), .C0(n5023), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_79_N3) );
  AOI2BB2X1 U6553 ( .B0(n389), .B1(K1[79]), .A0N(n5248), .A1N(n408), .Y(n5023)
         );
  XOR2X1 U6554 ( .A(n5249), .B(K1[13]), .Y(n5248) );
  CLKINVX1 U6555 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_79_), .Y(n5247) );
  CLKINVX1 U6556 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_94_), .Y(n5206) );
  OAI221X1 U6557 ( .A0(n330), .A1(n5210), .B0(n356), .B1(n5227), .C0(n5024), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_78_N3) );
  AOI2BB2X1 U6558 ( .B0(n389), .B1(K1[78]), .A0N(n5250), .A1N(n409), .Y(n5024)
         );
  XOR2X1 U6559 ( .A(n5251), .B(K1[12]), .Y(n5250) );
  CLKINVX1 U6560 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_78_), .Y(n5227) );
  OAI221X1 U6561 ( .A0(n330), .A1(n5213), .B0(n356), .B1(n5231), .C0(n5025), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_77_N3) );
  AOI2BB2X1 U6562 ( .B0(n389), .B1(K1[77]), .A0N(n5249), .A1N(n410), .Y(n5025)
         );
  XNOR2X1 U6563 ( .A(K1[11]), .B(n5252), .Y(n5249) );
  CLKINVX1 U6564 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_77_), .Y(n5231) );
  CLKINVX1 U6565 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_92_), .Y(n5213) );
  OAI221X1 U6566 ( .A0(n330), .A1(n5216), .B0(n356), .B1(n5235), .C0(n5026), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_76_N3) );
  AOI2BB2X1 U6567 ( .B0(n390), .B1(K1[76]), .A0N(n5251), .A1N(n408), .Y(n5026)
         );
  XNOR2X1 U6568 ( .A(K1[10]), .B(n5253), .Y(n5251) );
  CLKINVX1 U6569 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_76_), .Y(n5235) );
  CLKINVX1 U6570 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_91_), .Y(n5216) );
  OAI221X1 U6571 ( .A0(n331), .A1(n5218), .B0(n356), .B1(n5237), .C0(n5027), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_75_N3) );
  AOI22XL U6572 ( .A0(n5252), .A1(n414), .B0(n398), .B1(K1[75]), .Y(n5027) );
  XOR2X1 U6573 ( .A(K1[15]), .B(K1[9]), .Y(n5252) );
  CLKINVX1 U6574 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_75_), .Y(n5237) );
  CLKINVX1 U6575 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_90_), .Y(n5218) );
  OAI221X1 U6576 ( .A0(n331), .A1(n5224), .B0(n355), .B1(n5240), .C0(n5028), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_74_N3) );
  AOI22XL U6577 ( .A0(n5253), .A1(n414), .B0(n398), .B1(K1[74]), .Y(n5028) );
  XOR2X1 U6578 ( .A(K1[14]), .B(K1[8]), .Y(n5253) );
  CLKINVX1 U6579 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_74_), .Y(n5240) );
  CLKINVX1 U6580 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_89_), .Y(n5224) );
  OAI221X1 U6581 ( .A0(n331), .A1(n5226), .B0(n355), .B1(n5242), .C0(n5029), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_73_N3) );
  AOI22XL U6582 ( .A0(n414), .A1(K1[15]), .B0(n398), .B1(K1[73]), .Y(n5029) );
  CLKINVX1 U6583 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_73_), .Y(n5242) );
  CLKINVX1 U6584 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_88_), .Y(n5226) );
  OAI221X1 U6585 ( .A0(n5254), .A1(n341), .B0(n355), .B1(n5243), .C0(n5031), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_72_N3) );
  AOI22XL U6586 ( .A0(n414), .A1(K1[14]), .B0(n398), .B1(K1[72]), .Y(n5031) );
  CLKINVX1 U6587 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_72_), .Y(n5243) );
  XOR2X1 U6588 ( .A(n5210), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_95_), 
        .Y(n5254) );
  CLKINVX1 U6589 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_93_), .Y(n5210) );
  OAI221X1 U6590 ( .A0(n331), .A1(n5255), .B0(n355), .B1(n5256), .C0(n5034), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_71_N3) );
  AOI2BB2X1 U6591 ( .B0(n390), .B1(K1[71]), .A0N(n5257), .A1N(n409), .Y(n5034)
         );
  XOR2X1 U6592 ( .A(n5258), .B(K1[5]), .Y(n5257) );
  CLKINVX1 U6593 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_71_), .Y(n5256) );
  OAI221X1 U6594 ( .A0(n331), .A1(n5259), .B0(n355), .B1(n5260), .C0(n5037), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_70_N3) );
  AOI2BB2X1 U6595 ( .B0(n390), .B1(K1[70]), .A0N(n5261), .A1N(n410), .Y(n5037)
         );
  XOR2X1 U6596 ( .A(n5262), .B(K1[4]), .Y(n5261) );
  OAI221X1 U6597 ( .A0(n5263), .A1(n365), .B0(n5264), .B1(n345), .C0(n5040), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_7_N3) );
  AOI2BB2X1 U6598 ( .B0(n390), .B1(K1[7]), .A0N(n5265), .A1N(n408), .Y(n5040)
         );
  XOR2X1 U6599 ( .A(n4797), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_6_), 
        .Y(n5263) );
  OAI221X1 U6600 ( .A0(n331), .A1(n5266), .B0(n355), .B1(n5267), .C0(n5043), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_69_N3) );
  AOI2BB2X1 U6601 ( .B0(n390), .B1(K1[69]), .A0N(n5258), .A1N(n409), .Y(n5043)
         );
  XNOR2X1 U6602 ( .A(K1[3]), .B(n5268), .Y(n5258) );
  OAI221X1 U6603 ( .A0(n331), .A1(n5190), .B0(n355), .B1(n5269), .C0(n5045), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_68_N3) );
  AOI2BB2X1 U6604 ( .B0(n390), .B1(K1[68]), .A0N(n5262), .A1N(n410), .Y(n5045)
         );
  XNOR2X1 U6605 ( .A(K1[2]), .B(n5270), .Y(n5262) );
  CLKINVX1 U6606 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_99_), .Y(n5190) );
  OAI221X1 U6607 ( .A0(n331), .A1(n5194), .B0(n355), .B1(n5271), .C0(n5047), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_67_N3) );
  AOI22XL U6608 ( .A0(n5268), .A1(n414), .B0(n398), .B1(K1[67]), .Y(n5047) );
  XOR2X1 U6609 ( .A(K1[7]), .B(K1[1]), .Y(n5268) );
  CLKINVX1 U6610 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_98_), .Y(n5194) );
  OAI221X1 U6611 ( .A0(n331), .A1(n5197), .B0(n360), .B1(n5272), .C0(n5049), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_66_N3) );
  AOI22XL U6612 ( .A0(n5270), .A1(n414), .B0(n398), .B1(K1[66]), .Y(n5049) );
  XOR2X1 U6613 ( .A(K1[6]), .B(K1[0]), .Y(n5270) );
  CLKINVX1 U6614 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_97_), .Y(n5197) );
  OAI221X1 U6615 ( .A0(n331), .A1(n5199), .B0(n355), .B1(n5273), .C0(n5051), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_65_N3) );
  AOI22XL U6616 ( .A0(n414), .A1(K1[7]), .B0(n398), .B1(K1[65]), .Y(n5051) );
  CLKINVX1 U6617 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_96_), .Y(n5199) );
  OAI221X1 U6618 ( .A0(n5274), .A1(n341), .B0(n355), .B1(n5275), .C0(n5054), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_64_N3) );
  AOI22XL U6619 ( .A0(n414), .A1(K1[6]), .B0(n399), .B1(K1[64]), .Y(n5054) );
  XOR2X1 U6620 ( .A(n5259), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_103_), 
        .Y(n5274) );
  OAI221X1 U6621 ( .A0(n5276), .A1(n369), .B0(n5277), .B1(n345), .C0(n5056), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_63_N3) );
  AOI2BB2X1 U6622 ( .B0(n390), .B1(K1[63]), .A0N(n5278), .A1N(n408), .Y(n5056)
         );
  XOR2X1 U6623 ( .A(n4896), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_62_), 
        .Y(n5276) );
  OAI221X1 U6624 ( .A0(n5279), .A1(n341), .B0(n5280), .B1(n370), .C0(n5057), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_62_N3) );
  AOI2BB2X1 U6625 ( .B0(n390), .B1(K1[62]), .A0N(n5281), .A1N(n409), .Y(n5057)
         );
  XOR2X1 U6626 ( .A(n5282), .B(K1[109]), .Y(n5281) );
  OAI221X1 U6627 ( .A0(n5283), .A1(n341), .B0(n5284), .B1(n370), .C0(n5058), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_61_N3) );
  AOI2BB2X1 U6628 ( .B0(n390), .B1(K1[61]), .A0N(n5285), .A1N(n409), .Y(n5058)
         );
  XOR2X1 U6629 ( .A(n5278), .B(K1[110]), .Y(n5285) );
  XNOR2X1 U6630 ( .A(K1[108]), .B(n5286), .Y(n5278) );
  OAI221X1 U6631 ( .A0(n4659), .A1(n341), .B0(n5287), .B1(n369), .C0(n5059), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_60_N3) );
  AOI2BB2X1 U6632 ( .B0(n390), .B1(K1[60]), .A0N(n5282), .A1N(n408), .Y(n5059)
         );
  XNOR2X1 U6633 ( .A(K1[107]), .B(n5288), .Y(n5282) );
  OAI221X1 U6634 ( .A0(n5289), .A1(n342), .B0(n5290), .B1(n370), .C0(n5061), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_6_N3) );
  AOI2BB2X1 U6635 ( .B0(n390), .B1(K1[6]), .A0N(n5291), .A1N(n410), .Y(n5061)
         );
  XOR2X1 U6636 ( .A(n5292), .B(K1[117]), .Y(n5291) );
  OAI221X1 U6637 ( .A0(n5293), .A1(n342), .B0(n4856), .B1(n369), .C0(n5062), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_59_N3) );
  AOI2BB2X1 U6638 ( .B0(n390), .B1(K1[59]), .A0N(n5294), .A1N(n409), .Y(n5062)
         );
  XNOR2X1 U6639 ( .A(K1[110]), .B(n5286), .Y(n5294) );
  XOR2X1 U6640 ( .A(K1[104]), .B(K1[106]), .Y(n5286) );
  OAI221X1 U6641 ( .A0(n5295), .A1(n342), .B0(n5296), .B1(n370), .C0(n5063), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_58_N3) );
  AOI22XL U6642 ( .A0(n5288), .A1(n414), .B0(n398), .B1(K1[58]), .Y(n5063) );
  XOR2X1 U6643 ( .A(K1[111]), .B(K1[105]), .Y(n5288) );
  OAI221X1 U6644 ( .A0(n5297), .A1(n342), .B0(n5298), .B1(n370), .C0(n5065), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_57_N3) );
  AOI2BB2X1 U6645 ( .B0(n391), .B1(K1[57]), .A0N(n5299), .A1N(n409), .Y(n5065)
         );
  XNOR2X1 U6646 ( .A(K1[104]), .B(K1[110]), .Y(n5299) );
  OAI221X1 U6647 ( .A0(n5300), .A1(n342), .B0(n5301), .B1(n370), .C0(n5067), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_56_N3) );
  AOI22XL U6648 ( .A0(n414), .A1(K1[111]), .B0(n398), .B1(K1[56]), .Y(n5067)
         );
  OAI221X1 U6649 ( .A0(n5302), .A1(n369), .B0(n5290), .B1(n345), .C0(n5069), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_55_N3) );
  AOI2BB2X1 U6650 ( .B0(n391), .B1(K1[55]), .A0N(n5303), .A1N(n408), .Y(n5069)
         );
  CLKINVX1 U6651 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_7_), .Y(n5290)
         );
  XOR2X1 U6652 ( .A(n5300), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_54_), 
        .Y(n5302) );
  CLKINVX1 U6653 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_48_), .Y(n5300) );
  OAI221X1 U6654 ( .A0(n5304), .A1(n342), .B0(n5277), .B1(n370), .C0(n5070), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_54_N3) );
  AOI2BB2X1 U6655 ( .B0(n391), .B1(K1[54]), .A0N(n5305), .A1N(n410), .Y(n5070)
         );
  XOR2X1 U6656 ( .A(n5306), .B(K1[125]), .Y(n5305) );
  CLKINVX1 U6657 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_55_), .Y(n5277) );
  OAI221X1 U6658 ( .A0(n5307), .A1(n342), .B0(n5279), .B1(n370), .C0(n5071), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_53_N3) );
  AOI2BB2X1 U6659 ( .B0(n391), .B1(K1[53]), .A0N(n5308), .A1N(n410), .Y(n5071)
         );
  XOR2X1 U6660 ( .A(n5303), .B(K1[126]), .Y(n5308) );
  XNOR2X1 U6661 ( .A(K1[124]), .B(n5309), .Y(n5303) );
  CLKINVX1 U6662 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_54_), .Y(n5279) );
  OAI221X1 U6663 ( .A0(n4757), .A1(n342), .B0(n5283), .B1(n370), .C0(n5072), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_52_N3) );
  AOI2BB2X1 U6664 ( .B0(n391), .B1(K1[52]), .A0N(n5306), .A1N(n409), .Y(n5072)
         );
  XNOR2X1 U6665 ( .A(K1[123]), .B(n5310), .Y(n5306) );
  CLKINVX1 U6666 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_53_), .Y(n5283) );
  OAI221X1 U6667 ( .A0(n5311), .A1(n342), .B0(n4659), .B1(n370), .C0(n5073), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_51_N3) );
  AOI2BB2X1 U6668 ( .B0(n391), .B1(K1[51]), .A0N(n5312), .A1N(n408), .Y(n5073)
         );
  XNOR2X1 U6669 ( .A(K1[126]), .B(n5309), .Y(n5312) );
  XOR2X1 U6670 ( .A(K1[120]), .B(K1[122]), .Y(n5309) );
  CLKINVX1 U6671 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_52_), .Y(n4659) );
  OAI221X1 U6672 ( .A0(n5313), .A1(n342), .B0(n5293), .B1(n371), .C0(n5074), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_50_N3) );
  AOI22XL U6673 ( .A0(n5310), .A1(n414), .B0(n398), .B1(K1[50]), .Y(n5074) );
  XOR2X1 U6674 ( .A(K1[127]), .B(K1[121]), .Y(n5310) );
  CLKINVX1 U6675 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_51_), .Y(n5293) );
  OAI221X1 U6676 ( .A0(n5314), .A1(n342), .B0(n5304), .B1(n371), .C0(n5075), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_5_N3) );
  AOI2BB2X1 U6677 ( .B0(n391), .B1(K1[5]), .A0N(n5315), .A1N(n410), .Y(n5075)
         );
  XOR2X1 U6678 ( .A(n5265), .B(K1[118]), .Y(n5315) );
  XNOR2X1 U6679 ( .A(K1[116]), .B(n5316), .Y(n5265) );
  CLKINVX1 U6680 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_6_), .Y(n5304)
         );
  OAI221X1 U6681 ( .A0(n5317), .A1(n343), .B0(n5295), .B1(n370), .C0(n5077), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_49_N3) );
  AOI2BB2X1 U6682 ( .B0(n391), .B1(K1[49]), .A0N(n5318), .A1N(n408), .Y(n5077)
         );
  XNOR2X1 U6683 ( .A(K1[120]), .B(K1[126]), .Y(n5318) );
  CLKINVX1 U6684 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_50_), .Y(n5295) );
  OAI221X1 U6685 ( .A0(n4797), .A1(n343), .B0(n5297), .B1(n371), .C0(n5078), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_48_N3) );
  AOI22XL U6686 ( .A0(n414), .A1(K1[127]), .B0(n399), .B1(K1[48]), .Y(n5078)
         );
  CLKINVX1 U6687 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_49_), .Y(n5297) );
  CLKINVX1 U6688 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_0_), .Y(n4797)
         );
  OAI221X1 U6689 ( .A0(n5319), .A1(n369), .B0(n5280), .B1(n344), .C0(n5080), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_47_N3) );
  AOI2BB2X1 U6690 ( .B0(n391), .B1(K1[47]), .A0N(n5320), .A1N(n409), .Y(n5080)
         );
  CLKINVX1 U6691 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_63_), .Y(n5280) );
  XOR2X1 U6692 ( .A(n5321), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_46_), 
        .Y(n5319) );
  OAI221X1 U6693 ( .A0(n5284), .A1(n343), .B0(n5322), .B1(n371), .C0(n5082), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_46_N3) );
  AOI2BB2X1 U6694 ( .B0(n391), .B1(K1[46]), .A0N(n5323), .A1N(n408), .Y(n5082)
         );
  XOR2X1 U6695 ( .A(n5324), .B(K1[93]), .Y(n5323) );
  CLKINVX1 U6696 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_62_), .Y(n5284) );
  OAI221X1 U6697 ( .A0(n5287), .A1(n343), .B0(n5325), .B1(n371), .C0(n5084), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_45_N3) );
  AOI2BB2X1 U6698 ( .B0(n391), .B1(K1[45]), .A0N(n5326), .A1N(n410), .Y(n5084)
         );
  XOR2X1 U6699 ( .A(n5320), .B(K1[94]), .Y(n5326) );
  XNOR2X1 U6700 ( .A(K1[92]), .B(n5327), .Y(n5320) );
  CLKINVX1 U6701 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_61_), .Y(n5287) );
  OAI221X1 U6702 ( .A0(n4856), .A1(n343), .B0(n5328), .B1(n371), .C0(n5085), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_44_N3) );
  AOI2BB2X1 U6703 ( .B0(n391), .B1(K1[44]), .A0N(n5324), .A1N(n409), .Y(n5085)
         );
  XNOR2X1 U6704 ( .A(K1[91]), .B(n5329), .Y(n5324) );
  CLKINVX1 U6705 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_60_), .Y(n4856) );
  OAI221X1 U6706 ( .A0(n5296), .A1(n343), .B0(n5330), .B1(n371), .C0(n5086), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_43_N3) );
  AOI2BB2X1 U6707 ( .B0(n392), .B1(K1[43]), .A0N(n5331), .A1N(n409), .Y(n5086)
         );
  XNOR2X1 U6708 ( .A(K1[94]), .B(n5327), .Y(n5331) );
  XOR2X1 U6709 ( .A(K1[88]), .B(K1[90]), .Y(n5327) );
  CLKINVX1 U6710 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_59_), .Y(n5296) );
  OAI221X1 U6711 ( .A0(n5298), .A1(n343), .B0(n5332), .B1(n371), .C0(n5088), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_42_N3) );
  AOI22XL U6712 ( .A0(n5329), .A1(n414), .B0(n398), .B1(K1[42]), .Y(n5088) );
  XOR2X1 U6713 ( .A(K1[95]), .B(K1[89]), .Y(n5329) );
  CLKINVX1 U6714 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_58_), .Y(n5298) );
  OAI221X1 U6715 ( .A0(n5301), .A1(n343), .B0(n5333), .B1(n373), .C0(n5089), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_41_N3) );
  AOI2BB2X1 U6716 ( .B0(n392), .B1(K1[41]), .A0N(n5334), .A1N(n408), .Y(n5089)
         );
  XNOR2X1 U6717 ( .A(K1[88]), .B(K1[94]), .Y(n5334) );
  CLKINVX1 U6718 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_57_), .Y(n5301) );
  OAI221X1 U6719 ( .A0(n4896), .A1(n343), .B0(n5335), .B1(n371), .C0(n5090), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_40_N3) );
  AOI22XL U6720 ( .A0(n414), .A1(K1[95]), .B0(n398), .B1(K1[40]), .Y(n5090) );
  CLKINVX1 U6721 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_56_), .Y(n4896) );
  OAI221X1 U6722 ( .A0(n5336), .A1(n343), .B0(n5307), .B1(n371), .C0(n5091), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_4_N3) );
  AOI2BB2X1 U6723 ( .B0(n392), .B1(K1[4]), .A0N(n5292), .A1N(n410), .Y(n5091)
         );
  XNOR2X1 U6724 ( .A(K1[115]), .B(n5337), .Y(n5292) );
  CLKINVX1 U6725 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_5_), .Y(n5307)
         );
  OAI221X1 U6726 ( .A0(n5338), .A1(n369), .B0(n5339), .B1(n345), .C0(n5094), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_39_N3) );
  AOI2BB2X1 U6727 ( .B0(n392), .B1(K1[39]), .A0N(n5340), .A1N(n410), .Y(n5094)
         );
  XOR2X1 U6728 ( .A(n5341), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_38_), 
        .Y(n5338) );
  OAI221X1 U6729 ( .A0(n5342), .A1(n342), .B0(n5264), .B1(n371), .C0(n5095), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_38_N3) );
  AOI2BB2X1 U6730 ( .B0(n392), .B1(K1[38]), .A0N(n5343), .A1N(n408), .Y(n5095)
         );
  XOR2X1 U6731 ( .A(n5344), .B(K1[69]), .Y(n5343) );
  CLKINVX1 U6732 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_39_), .Y(n5264) );
  OAI221X1 U6733 ( .A0(n5345), .A1(n342), .B0(n5289), .B1(n371), .C0(n5096), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_37_N3) );
  AOI2BB2X1 U6734 ( .B0(n392), .B1(K1[37]), .A0N(n5346), .A1N(n410), .Y(n5096)
         );
  XOR2X1 U6735 ( .A(n5340), .B(K1[70]), .Y(n5346) );
  XNOR2X1 U6736 ( .A(K1[68]), .B(n5347), .Y(n5340) );
  CLKINVX1 U6737 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_38_), .Y(n5289) );
  OAI221X1 U6738 ( .A0(n5348), .A1(n344), .B0(n5314), .B1(n372), .C0(n5097), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_36_N3) );
  AOI2BB2X1 U6739 ( .B0(n392), .B1(K1[36]), .A0N(n5344), .A1N(n410), .Y(n5097)
         );
  XNOR2X1 U6740 ( .A(K1[67]), .B(n5349), .Y(n5344) );
  CLKINVX1 U6741 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_37_), .Y(n5314) );
  OAI221X1 U6742 ( .A0(n5350), .A1(n343), .B0(n5336), .B1(n372), .C0(n5099), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_35_N3) );
  AOI2BB2X1 U6743 ( .B0(n392), .B1(K1[35]), .A0N(n5351), .A1N(n410), .Y(n5099)
         );
  XNOR2X1 U6744 ( .A(K1[70]), .B(n5347), .Y(n5351) );
  XOR2X1 U6745 ( .A(K1[64]), .B(K1[66]), .Y(n5347) );
  CLKINVX1 U6746 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_36_), .Y(n5336) );
  OAI221X1 U6747 ( .A0(n5352), .A1(n344), .B0(n5353), .B1(n372), .C0(n5101), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_34_N3) );
  AOI22XL U6748 ( .A0(n5349), .A1(n414), .B0(n398), .B1(K1[34]), .Y(n5101) );
  XOR2X1 U6749 ( .A(K1[71]), .B(K1[65]), .Y(n5349) );
  OAI221X1 U6750 ( .A0(n5354), .A1(n344), .B0(n5355), .B1(n374), .C0(n5103), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_33_N3) );
  AOI2BB2X1 U6751 ( .B0(n392), .B1(K1[33]), .A0N(n5356), .A1N(n409), .Y(n5103)
         );
  XNOR2X1 U6752 ( .A(K1[64]), .B(K1[70]), .Y(n5356) );
  OAI221X1 U6753 ( .A0(n5357), .A1(n343), .B0(n5358), .B1(n374), .C0(n5104), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_32_N3) );
  AOI22XL U6754 ( .A0(n414), .A1(K1[71]), .B0(n397), .B1(K1[32]), .Y(n5104) );
  OAI221X1 U6755 ( .A0(n5359), .A1(n369), .B0(n5322), .B1(n345), .C0(n5106), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_31_N3) );
  AOI2BB2X1 U6756 ( .B0(n392), .B1(K1[31]), .A0N(n5360), .A1N(n408), .Y(n5106)
         );
  CLKINVX1 U6757 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_47_), .Y(n5322) );
  XOR2X1 U6758 ( .A(n5245), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_30_), 
        .Y(n5359) );
  CLKINVX1 U6759 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_24_), .Y(n5245) );
  OAI221X1 U6760 ( .A0(n5325), .A1(n344), .B0(n5361), .B1(n376), .C0(n5108), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_30_N3) );
  AOI2BB2X1 U6761 ( .B0(n395), .B1(K1[30]), .A0N(n5362), .A1N(n408), .Y(n5108)
         );
  XOR2X1 U6762 ( .A(n5363), .B(K1[77]), .Y(n5362) );
  CLKINVX1 U6763 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_46_), .Y(n5325) );
  OAI221X1 U6764 ( .A0(n5353), .A1(n344), .B0(n4757), .B1(n376), .C0(n5109), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_3_N3) );
  AOI2BB2X1 U6765 ( .B0(n392), .B1(K1[3]), .A0N(n5364), .A1N(n410), .Y(n5109)
         );
  XNOR2X1 U6766 ( .A(K1[118]), .B(n5316), .Y(n5364) );
  XOR2X1 U6767 ( .A(K1[112]), .B(K1[114]), .Y(n5316) );
  CLKINVX1 U6768 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_4_), .Y(n4757)
         );
  CLKINVX1 U6769 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_35_), .Y(n5353) );
  OAI221X1 U6770 ( .A0(n5328), .A1(n344), .B0(n5365), .B1(n377), .C0(n5111), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_29_N3) );
  AOI2BB2X1 U6771 ( .B0(n392), .B1(K1[29]), .A0N(n5366), .A1N(n408), .Y(n5111)
         );
  XOR2X1 U6772 ( .A(n5360), .B(K1[78]), .Y(n5366) );
  XNOR2X1 U6773 ( .A(K1[76]), .B(n5367), .Y(n5360) );
  CLKINVX1 U6774 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_45_), .Y(n5328) );
  OAI221X1 U6775 ( .A0(n5330), .A1(n344), .B0(n5368), .B1(n369), .C0(n5112), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_28_N3) );
  AOI2BB2X1 U6776 ( .B0(n393), .B1(K1[28]), .A0N(n5363), .A1N(n409), .Y(n5112)
         );
  XNOR2X1 U6777 ( .A(K1[75]), .B(n5369), .Y(n5363) );
  CLKINVX1 U6778 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_44_), .Y(n5330) );
  OAI221X1 U6779 ( .A0(n5332), .A1(n344), .B0(n5370), .B1(n377), .C0(n5113), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_27_N3) );
  AOI2BB2X1 U6780 ( .B0(n393), .B1(K1[27]), .A0N(n5371), .A1N(n410), .Y(n5113)
         );
  XNOR2X1 U6781 ( .A(K1[78]), .B(n5367), .Y(n5371) );
  XOR2X1 U6782 ( .A(K1[72]), .B(K1[74]), .Y(n5367) );
  CLKINVX1 U6783 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_43_), .Y(n5332) );
  OAI221X1 U6784 ( .A0(n5333), .A1(n325), .B0(n5372), .B1(n377), .C0(n5115), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_26_N3) );
  AOI22XL U6785 ( .A0(n5369), .A1(n414), .B0(n397), .B1(K1[26]), .Y(n5115) );
  XOR2X1 U6786 ( .A(K1[79]), .B(K1[73]), .Y(n5369) );
  CLKINVX1 U6787 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_42_), .Y(n5333) );
  OAI221X1 U6788 ( .A0(n5335), .A1(n343), .B0(n5373), .B1(n377), .C0(n5116), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_25_N3) );
  AOI2BB2X1 U6789 ( .B0(n393), .B1(K1[25]), .A0N(n5374), .A1N(n408), .Y(n5116)
         );
  XNOR2X1 U6790 ( .A(K1[72]), .B(K1[78]), .Y(n5374) );
  CLKINVX1 U6791 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_41_), .Y(n5335) );
  OAI221X1 U6792 ( .A0(n5321), .A1(n327), .B0(n5219), .B1(n377), .C0(n5117), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_24_N3) );
  AOI22XL U6793 ( .A0(n414), .A1(K1[79]), .B0(n397), .B1(K1[24]), .Y(n5117) );
  CLKINVX1 U6794 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_25_), .Y(n5219) );
  CLKINVX1 U6795 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_40_), .Y(n5321) );
  OAI221X1 U6796 ( .A0(n5375), .A1(n369), .B0(n5376), .B1(n345), .C0(n5120), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_23_N3) );
  AOI2BB2X1 U6797 ( .B0(n393), .B1(K1[23]), .A0N(n5377), .A1N(n410), .Y(n5120)
         );
  XOR2X1 U6798 ( .A(n5357), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_22_), 
        .Y(n5375) );
  CLKINVX1 U6799 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_16_), .Y(n5357) );
  OAI221X1 U6800 ( .A0(n5378), .A1(n344), .B0(n5339), .B1(n377), .C0(n5122), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_22_N3) );
  AOI2BB2X1 U6801 ( .B0(n393), .B1(K1[22]), .A0N(n5379), .A1N(n409), .Y(n5122)
         );
  XOR2X1 U6802 ( .A(n5380), .B(K1[101]), .Y(n5379) );
  CLKINVX1 U6803 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_23_), .Y(n5339) );
  OAI221X1 U6804 ( .A0(n5381), .A1(n333), .B0(n5342), .B1(n377), .C0(n5123), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_21_N3) );
  AOI2BB2X1 U6805 ( .B0(n393), .B1(K1[21]), .A0N(n5382), .A1N(n409), .Y(n5123)
         );
  XOR2X1 U6806 ( .A(n5377), .B(K1[102]), .Y(n5382) );
  XNOR2X1 U6807 ( .A(K1[100]), .B(n5383), .Y(n5377) );
  CLKINVX1 U6808 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_22_), .Y(n5342) );
  OAI221X1 U6809 ( .A0(n5384), .A1(n344), .B0(n5345), .B1(n377), .C0(n5124), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_20_N3) );
  AOI2BB2X1 U6810 ( .B0(n393), .B1(K1[20]), .A0N(n5380), .A1N(n409), .Y(n5124)
         );
  XNOR2X1 U6811 ( .A(K1[99]), .B(n5385), .Y(n5380) );
  CLKINVX1 U6812 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_21_), .Y(n5345) );
  OAI221X1 U6813 ( .A0(n5355), .A1(n344), .B0(n5311), .B1(n377), .C0(n5125), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_2_N3) );
  AOI22XL U6814 ( .A0(n5337), .A1(n414), .B0(n397), .B1(K1[2]), .Y(n5125) );
  XOR2X1 U6815 ( .A(K1[119]), .B(K1[113]), .Y(n5337) );
  CLKINVX1 U6816 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_3_), .Y(n5311)
         );
  CLKINVX1 U6817 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_34_), .Y(n5355) );
  OAI221X1 U6818 ( .A0(n5386), .A1(n328), .B0(n5348), .B1(n377), .C0(n5127), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_19_N3) );
  AOI2BB2X1 U6819 ( .B0(n393), .B1(K1[19]), .A0N(n5387), .A1N(n408), .Y(n5127)
         );
  XNOR2X1 U6820 ( .A(K1[102]), .B(n5383), .Y(n5387) );
  XOR2X1 U6821 ( .A(K1[96]), .B(K1[98]), .Y(n5383) );
  CLKINVX1 U6822 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_20_), .Y(n5348) );
  OAI221X1 U6823 ( .A0(n5220), .A1(n344), .B0(n5350), .B1(n377), .C0(n5128), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_18_N3) );
  AOI22XL U6824 ( .A0(n5385), .A1(n414), .B0(n397), .B1(K1[18]), .Y(n5128) );
  XOR2X1 U6825 ( .A(K1[103]), .B(K1[97]), .Y(n5385) );
  CLKINVX1 U6826 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_19_), .Y(n5350) );
  CLKINVX1 U6827 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_10_), .Y(n5220) );
  OAI221X1 U6828 ( .A0(n5246), .A1(n326), .B0(n5352), .B1(n376), .C0(n5129), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_17_N3) );
  AOI2BB2X1 U6829 ( .B0(n393), .B1(K1[17]), .A0N(n5388), .A1N(n410), .Y(n5129)
         );
  XNOR2X1 U6830 ( .A(K1[96]), .B(K1[102]), .Y(n5388) );
  CLKINVX1 U6831 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_18_), .Y(n5352) );
  CLKINVX1 U6832 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_9_), .Y(n5246)
         );
  OAI221X1 U6833 ( .A0(n5389), .A1(n332), .B0(n5354), .B1(n376), .C0(n5130), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_16_N3) );
  AOI22XL U6834 ( .A0(n414), .A1(K1[103]), .B0(n397), .B1(K1[16]), .Y(n5130)
         );
  CLKINVX1 U6835 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_17_), .Y(n5354) );
  OAI221X1 U6836 ( .A0(n5390), .A1(n369), .B0(n5361), .B1(n345), .C0(n5132), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_15_N3) );
  AOI2BB2X1 U6837 ( .B0(n393), .B1(K1[15]), .A0N(n5391), .A1N(n410), .Y(n5132)
         );
  CLKINVX1 U6838 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_31_), .Y(n5361) );
  XOR2X1 U6839 ( .A(n5389), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_14_), 
        .Y(n5390) );
  CLKINVX1 U6840 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_8_), .Y(n5389)
         );
  OAI221X1 U6841 ( .A0(n5365), .A1(n340), .B0(n5376), .B1(n376), .C0(n5133), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_14_N3) );
  AOI2BB2X1 U6842 ( .B0(n393), .B1(K1[14]), .A0N(n5392), .A1N(n409), .Y(n5133)
         );
  XOR2X1 U6843 ( .A(n5393), .B(K1[85]), .Y(n5392) );
  CLKINVX1 U6844 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_15_), .Y(n5376) );
  CLKINVX1 U6845 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_30_), .Y(n5365) );
  OAI221X1 U6846 ( .A0(n5368), .A1(n335), .B0(n5378), .B1(n376), .C0(n5134), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_13_N3) );
  AOI2BB2X1 U6847 ( .B0(n393), .B1(K1[13]), .A0N(n5394), .A1N(n409), .Y(n5134)
         );
  XOR2X1 U6848 ( .A(n5391), .B(K1[86]), .Y(n5394) );
  XNOR2X1 U6849 ( .A(K1[84]), .B(n5395), .Y(n5391) );
  CLKINVX1 U6850 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_14_), .Y(n5378) );
  CLKINVX1 U6851 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_29_), .Y(n5368) );
  OAI221X1 U6852 ( .A0(n335), .A1(n5396), .B0(n359), .B1(n5397), .C0(n5137), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_127_N3) );
  AOI2BB2X1 U6853 ( .B0(n394), .B1(K1[127]), .A0N(n5398), .A1N(n408), .Y(n5137) );
  XOR2X1 U6854 ( .A(n5399), .B(K1[61]), .Y(n5398) );
  CLKINVX1 U6855 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_127_), .Y(
        n5397) );
  OAI221X1 U6856 ( .A0(n335), .A1(n5400), .B0(n359), .B1(n5401), .C0(n5140), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_126_N3) );
  AOI2BB2X1 U6857 ( .B0(n394), .B1(K1[126]), .A0N(n5402), .A1N(n410), .Y(n5140) );
  XOR2X1 U6858 ( .A(n5403), .B(K1[60]), .Y(n5402) );
  OAI221X1 U6859 ( .A0(n336), .A1(n5404), .B0(n359), .B1(n5405), .C0(n5143), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_125_N3) );
  AOI2BB2X1 U6860 ( .B0(n394), .B1(K1[125]), .A0N(n5399), .A1N(n408), .Y(n5143) );
  XNOR2X1 U6861 ( .A(K1[59]), .B(n5406), .Y(n5399) );
  OAI221X1 U6862 ( .A0(n336), .A1(n5407), .B0(n359), .B1(n5408), .C0(n5146), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_124_N3) );
  AOI2BB2X1 U6863 ( .B0(n394), .B1(K1[124]), .A0N(n5403), .A1N(n409), .Y(n5146) );
  XNOR2X1 U6864 ( .A(K1[58]), .B(n5409), .Y(n5403) );
  OAI221X1 U6865 ( .A0(n332), .A1(n5410), .B0(n359), .B1(n5411), .C0(n5149), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_123_N3) );
  AOI22XL U6866 ( .A0(n5406), .A1(n414), .B0(n397), .B1(K1[123]), .Y(n5149) );
  XOR2X1 U6867 ( .A(K1[63]), .B(K1[57]), .Y(n5406) );
  OAI221X1 U6868 ( .A0(n335), .A1(n5412), .B0(n360), .B1(n5413), .C0(n5152), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_122_N3) );
  AOI22XL U6869 ( .A0(n5409), .A1(n414), .B0(n396), .B1(K1[122]), .Y(n5152) );
  XOR2X1 U6870 ( .A(K1[62]), .B(K1[56]), .Y(n5409) );
  OAI221X1 U6871 ( .A0(n335), .A1(n5414), .B0(n360), .B1(n5415), .C0(n5155), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_121_N3) );
  AOI22XL U6872 ( .A0(n414), .A1(K1[63]), .B0(n397), .B1(K1[121]), .Y(n5155)
         );
  OAI221X1 U6873 ( .A0(n5416), .A1(n331), .B0(n360), .B1(n5417), .C0(n5158), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_120_N3) );
  AOI22XL U6874 ( .A0(n414), .A1(K1[62]), .B0(n396), .B1(K1[120]), .Y(n5158)
         );
  XOR2X1 U6875 ( .A(n5400), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_119_), 
        .Y(n5416) );
  OAI221X1 U6876 ( .A0(n5370), .A1(n330), .B0(n5381), .B1(n376), .C0(n5159), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_12_N3) );
  AOI2BB2X1 U6877 ( .B0(n394), .B1(K1[12]), .A0N(n5393), .A1N(n410), .Y(n5159)
         );
  XNOR2X1 U6878 ( .A(K1[83]), .B(n5418), .Y(n5393) );
  CLKINVX1 U6879 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_13_), .Y(n5381) );
  CLKINVX1 U6880 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_28_), .Y(n5370) );
  OAI221X1 U6881 ( .A0(n334), .A1(n5260), .B0(n360), .B1(n5419), .C0(n5161), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_119_N3) );
  AOI2BB2X1 U6882 ( .B0(n394), .B1(K1[119]), .A0N(n5420), .A1N(n410), .Y(n5161) );
  XOR2X1 U6883 ( .A(n5421), .B(K1[53]), .Y(n5420) );
  CLKINVX1 U6884 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_119_), .Y(
        n5419) );
  CLKINVX1 U6885 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_70_), .Y(n5260) );
  OAI221X1 U6886 ( .A0(n335), .A1(n5267), .B0(n360), .B1(n5396), .C0(n5162), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_118_N3) );
  AOI2BB2X1 U6887 ( .B0(n394), .B1(K1[118]), .A0N(n5422), .A1N(n409), .Y(n5162) );
  XOR2X1 U6888 ( .A(n5423), .B(K1[52]), .Y(n5422) );
  CLKINVX1 U6889 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_118_), .Y(
        n5396) );
  OAI221X1 U6890 ( .A0(n335), .A1(n5269), .B0(n360), .B1(n5400), .C0(n5163), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_117_N3) );
  AOI2BB2X1 U6891 ( .B0(n394), .B1(K1[117]), .A0N(n5421), .A1N(n408), .Y(n5163) );
  XNOR2X1 U6892 ( .A(K1[51]), .B(n5424), .Y(n5421) );
  CLKINVX1 U6893 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_117_), .Y(
        n5400) );
  CLKINVX1 U6894 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_68_), .Y(n5269) );
  OAI221X1 U6895 ( .A0(n334), .A1(n5271), .B0(n360), .B1(n5404), .C0(n5164), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_116_N3) );
  AOI2BB2X1 U6896 ( .B0(n394), .B1(K1[116]), .A0N(n5423), .A1N(n408), .Y(n5164) );
  XNOR2X1 U6897 ( .A(K1[50]), .B(n5425), .Y(n5423) );
  CLKINVX1 U6898 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_116_), .Y(
        n5404) );
  CLKINVX1 U6899 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_67_), .Y(n5271) );
  OAI221X1 U6900 ( .A0(n334), .A1(n5272), .B0(n360), .B1(n5407), .C0(n5165), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_115_N3) );
  AOI22XL U6901 ( .A0(n5424), .A1(n414), .B0(n396), .B1(K1[115]), .Y(n5165) );
  XOR2X1 U6902 ( .A(K1[55]), .B(K1[49]), .Y(n5424) );
  CLKINVX1 U6903 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_115_), .Y(
        n5407) );
  CLKINVX1 U6904 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_66_), .Y(n5272) );
  OAI221X1 U6905 ( .A0(n334), .A1(n5273), .B0(n360), .B1(n5410), .C0(n5166), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_114_N3) );
  AOI22XL U6906 ( .A0(n5425), .A1(n414), .B0(n397), .B1(K1[114]), .Y(n5166) );
  XOR2X1 U6907 ( .A(K1[54]), .B(K1[48]), .Y(n5425) );
  CLKINVX1 U6908 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_114_), .Y(
        n5410) );
  CLKINVX1 U6909 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_65_), .Y(n5273) );
  OAI221X1 U6910 ( .A0(n333), .A1(n5275), .B0(n360), .B1(n5412), .C0(n5167), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_113_N3) );
  AOI22XL U6911 ( .A0(n414), .A1(K1[55]), .B0(n396), .B1(K1[113]), .Y(n5167)
         );
  CLKINVX1 U6912 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_113_), .Y(
        n5412) );
  CLKINVX1 U6913 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_64_), .Y(n5275) );
  OAI221X1 U6914 ( .A0(n5426), .A1(n334), .B0(n360), .B1(n5414), .C0(n5169), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_112_N3) );
  AOI22XL U6915 ( .A0(n414), .A1(K1[54]), .B0(n396), .B1(K1[112]), .Y(n5169)
         );
  CLKINVX1 U6916 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_112_), .Y(
        n5414) );
  XOR2X1 U6917 ( .A(n5267), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_71_), 
        .Y(n5426) );
  CLKINVX1 U6918 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_69_), .Y(n5267) );
  OAI221X1 U6919 ( .A0(n334), .A1(n5401), .B0(n361), .B1(n5427), .C0(n5171), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_111_N3) );
  AOI2BB2X1 U6920 ( .B0(n394), .B1(K1[111]), .A0N(n5428), .A1N(n408), .Y(n5171) );
  XOR2X1 U6921 ( .A(n5429), .B(K1[45]), .Y(n5428) );
  CLKINVX1 U6922 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_111_), .Y(
        n5427) );
  CLKINVX1 U6923 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_126_), .Y(
        n5401) );
  OAI221X1 U6924 ( .A0(n333), .A1(n5405), .B0(n361), .B1(n5201), .C0(n5172), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_110_N3) );
  AOI2BB2X1 U6925 ( .B0(n394), .B1(K1[110]), .A0N(n5430), .A1N(n410), .Y(n5172) );
  XOR2X1 U6926 ( .A(n5431), .B(K1[44]), .Y(n5430) );
  CLKINVX1 U6927 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_110_), .Y(
        n5201) );
  OAI221X1 U6928 ( .A0(n5372), .A1(n344), .B0(n5384), .B1(n376), .C0(n5173), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_11_N3) );
  AOI2BB2X1 U6929 ( .B0(n394), .B1(K1[11]), .A0N(n5432), .A1N(n408), .Y(n5173)
         );
  XOR2X1 U6930 ( .A(n5222), .B(n5395), .Y(n5432) );
  XOR2X1 U6931 ( .A(K1[80]), .B(K1[82]), .Y(n5395) );
  CLKINVX1 U6932 ( .A(K1[86]), .Y(n5222) );
  CLKINVX1 U6933 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_12_), .Y(n5384) );
  CLKINVX1 U6934 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_27_), .Y(n5372) );
  OAI221X1 U6935 ( .A0(n333), .A1(n5408), .B0(n361), .B1(n5205), .C0(n5174), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_109_N3) );
  AOI2BB2X1 U6936 ( .B0(n395), .B1(K1[109]), .A0N(n5429), .A1N(n409), .Y(n5174) );
  XNOR2X1 U6937 ( .A(K1[43]), .B(n5433), .Y(n5429) );
  CLKINVX1 U6938 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_109_), .Y(
        n5205) );
  CLKINVX1 U6939 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_124_), .Y(
        n5408) );
  OAI221X1 U6940 ( .A0(n333), .A1(n5411), .B0(n361), .B1(n5209), .C0(n5175), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_108_N3) );
  AOI2BB2X1 U6941 ( .B0(n395), .B1(K1[108]), .A0N(n5431), .A1N(n408), .Y(n5175) );
  XNOR2X1 U6942 ( .A(K1[42]), .B(n5434), .Y(n5431) );
  CLKINVX1 U6943 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_108_), .Y(
        n5209) );
  CLKINVX1 U6944 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_123_), .Y(
        n5411) );
  OAI221X1 U6945 ( .A0(n333), .A1(n5413), .B0(n361), .B1(n5212), .C0(n5176), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_107_N3) );
  AOI22XL U6946 ( .A0(n5433), .A1(n414), .B0(n396), .B1(K1[107]), .Y(n5176) );
  XOR2X1 U6947 ( .A(K1[47]), .B(K1[41]), .Y(n5433) );
  CLKINVX1 U6948 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_107_), .Y(
        n5212) );
  CLKINVX1 U6949 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_122_), .Y(
        n5413) );
  OAI221X1 U6950 ( .A0(n333), .A1(n5415), .B0(n361), .B1(n5215), .C0(n5177), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_106_N3) );
  AOI22XL U6951 ( .A0(n5434), .A1(n414), .B0(n396), .B1(K1[106]), .Y(n5177) );
  XOR2X1 U6952 ( .A(K1[46]), .B(K1[40]), .Y(n5434) );
  CLKINVX1 U6953 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_106_), .Y(
        n5215) );
  CLKINVX1 U6954 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_121_), .Y(
        n5415) );
  OAI221X1 U6955 ( .A0(n333), .A1(n5417), .B0(n361), .B1(n5217), .C0(n5178), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_105_N3) );
  AOI22XL U6956 ( .A0(n414), .A1(K1[47]), .B0(n396), .B1(K1[105]), .Y(n5178)
         );
  CLKINVX1 U6957 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_105_), .Y(
        n5217) );
  CLKINVX1 U6958 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_120_), .Y(
        n5417) );
  OAI221X1 U6959 ( .A0(n5435), .A1(n336), .B0(n361), .B1(n5223), .C0(n5180), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_104_N3) );
  AOI22XL U6960 ( .A0(n414), .A1(K1[46]), .B0(n396), .B1(K1[104]), .Y(n5180)
         );
  CLKINVX1 U6961 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_104_), .Y(
        n5223) );
  XOR2X1 U6962 ( .A(n5405), .B(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_127_), 
        .Y(n5435) );
  CLKINVX1 U6963 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_125_), .Y(
        n5405) );
  OAI221X1 U6964 ( .A0(n333), .A1(n5232), .B0(n361), .B1(n5436), .C0(n5182), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_103_N3) );
  AOI2BB2X1 U6965 ( .B0(n395), .B1(K1[103]), .A0N(n5437), .A1N(n409), .Y(n5182) );
  XOR2X1 U6966 ( .A(n5438), .B(K1[37]), .Y(n5437) );
  CLKINVX1 U6967 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_103_), .Y(
        n5436) );
  CLKINVX1 U6968 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_86_), .Y(n5232) );
  OAI221X1 U6969 ( .A0(n333), .A1(n5200), .B0(n361), .B1(n5255), .C0(n5183), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_102_N3) );
  AOI2BB2X1 U6970 ( .B0(n395), .B1(K1[102]), .A0N(n5439), .A1N(n408), .Y(n5183) );
  XOR2X1 U6971 ( .A(n5440), .B(K1[36]), .Y(n5439) );
  CLKINVX1 U6972 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_102_), .Y(
        n5255) );
  CLKINVX1 U6973 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_85_), .Y(n5200) );
  OAI221X1 U6974 ( .A0(n333), .A1(n5238), .B0(n361), .B1(n5259), .C0(n5184), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_101_N3) );
  AOI2BB2X1 U6975 ( .B0(n395), .B1(K1[101]), .A0N(n5438), .A1N(n410), .Y(n5184) );
  XNOR2X1 U6976 ( .A(K1[35]), .B(n5191), .Y(n5438) );
  XOR2X1 U6977 ( .A(K1[39]), .B(K1[33]), .Y(n5191) );
  CLKINVX1 U6978 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_101_), .Y(
        n5259) );
  CLKINVX1 U6979 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_84_), .Y(n5238) );
  OAI221X1 U6980 ( .A0(n333), .A1(n5241), .B0(n361), .B1(n5266), .C0(n5185), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_100_N3) );
  AOI2BB2X1 U6981 ( .B0(n395), .B1(K1[100]), .A0N(n5440), .A1N(n409), .Y(n5185) );
  XNOR2X1 U6982 ( .A(K1[34]), .B(n5195), .Y(n5440) );
  XOR2X1 U6983 ( .A(K1[38]), .B(K1[32]), .Y(n5195) );
  CLKINVX1 U6984 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_100_), .Y(
        n5266) );
  CLKINVX1 U6985 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_83_), .Y(n5241) );
  OAI221X1 U6986 ( .A0(n5373), .A1(n329), .B0(n5386), .B1(n376), .C0(n5186), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_10_N3) );
  AOI22XL U6987 ( .A0(n5418), .A1(n414), .B0(n396), .B1(K1[10]), .Y(n5186) );
  XOR2X1 U6988 ( .A(K1[87]), .B(K1[81]), .Y(n5418) );
  CLKINVX1 U6989 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_11_), .Y(n5386) );
  CLKINVX1 U6990 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_26_), .Y(n5373) );
  OAI221X1 U6991 ( .A0(n5358), .A1(n340), .B0(n5313), .B1(n376), .C0(n5187), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_1_N3) );
  AOI2BB2X1 U6992 ( .B0(n395), .B1(K1[1]), .A0N(n5441), .A1N(n408), .Y(n5187)
         );
  XNOR2X1 U6993 ( .A(K1[112]), .B(K1[118]), .Y(n5441) );
  CLKINVX1 U6994 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_2_), .Y(n5313)
         );
  CLKINVX1 U6995 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_33_), .Y(n5358) );
  OAI221X1 U6996 ( .A0(n5341), .A1(n345), .B0(n5317), .B1(n376), .C0(n5188), 
        .Y(Inst_forkAE_CipherInst_KE_RS2_1_SFF_0_N3) );
  AOI22XL U6997 ( .A0(n414), .A1(K1[119]), .B0(n396), .B1(K1[0]), .Y(n5188) );
  CLKINVX1 U6998 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_1_), .Y(n5317)
         );
  CLKINVX1 U6999 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM2_1_Inv_32_), .Y(n5341) );
  CLKINVX1 U7000 ( .A(n5442), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_99_N3) );
  AOI222XL U7001 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[99]), .B0(n347), .B1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[83]), .C0(n414), .C1(
        N[35]), .Y(n5442) );
  CLKINVX1 U7002 ( .A(n5444), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_98_N3) );
  AOI221XL U7003 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[98]), .B0(n411), .B1(N[34]), .C0(n5445), .Y(n5444) );
  CLKINVX1 U7004 ( .A(n5446), .Y(n5445) );
  AOI32XL U7005 ( .A0(n395), .A1(n4958), .A2(n1998), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[82]), .B1(n354), .Y(n5446) );
  NOR3X1 U7006 ( .A(dec), .B(enc), .C(n1986), .Y(n1998) );
  NOR2BX1 U7007 ( .AN(gen_tag), .B(a_data), .Y(n4958) );
  CLKINVX1 U7008 ( .A(n5447), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_97_N3) );
  AOI221XL U7009 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[97]), .B0(n412), .B1(N[33]), .C0(n5448), .Y(n5447) );
  OAI32XL U7010 ( .A0(n1986), .A1(n1972), .A2(n5449), .B0(n5450), .B1(n342), 
        .Y(n5448) );
  CLKINVX1 U7011 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[81]), .Y(n5450)
         );
  CLKINVX1 U7012 ( .A(a_data), .Y(n1972) );
  CLKINVX1 U7013 ( .A(n5451), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_96_N3) );
  AOI221XL U7014 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[96]), .B0(n413), .B1(N[32]), .C0(n5452), .Y(n5451) );
  OAI32XL U7015 ( .A0(n5453), .A1(n255), .A2(n1986), .B0(n5454), .B1(n341), 
        .Y(n5452) );
  CLKINVX1 U7016 ( .A(Inst_forkAE_ControlInst_fsm_state_0_), .Y(n1986) );
  AOI21X1 U7017 ( .A0(n145), .A1(n1982), .B0(n180), .Y(n5453) );
  OR3X1 U7018 ( .A(enc), .B(gen_tag), .C(dec), .Y(n1982) );
  CLKINVX1 U7019 ( .A(n5455), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_95_N3) );
  AOI221XL U7020 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[95]), .B0(n413), .B1(N[31]), .C0(n5456), .Y(n5455) );
  OAI2B2X1 U7021 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[111]), .A0(
        n325), .B0(n5457), .B1(n5449), .Y(n5456) );
  CLKINVX1 U7022 ( .A(n5458), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_94_N3) );
  AOI221XL U7023 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[94]), .B0(n413), .B1(N[30]), .C0(n5459), .Y(n5458) );
  OAI2B2X1 U7024 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[110]), .A0(
        n325), .B0(n5460), .B1(n5449), .Y(n5459) );
  CLKINVX1 U7025 ( .A(n5461), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_93_N3) );
  AOI221XL U7026 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[93]), .B0(n413), .B1(N[29]), .C0(n5462), .Y(n5461) );
  OAI2B2X1 U7027 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[109]), .A0(
        n326), .B0(n5463), .B1(n5449), .Y(n5462) );
  CLKINVX1 U7028 ( .A(n5464), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_92_N3) );
  AOI221XL U7029 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[92]), .B0(n413), .B1(N[28]), .C0(n5465), .Y(n5464) );
  OAI2B2X1 U7030 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[108]), .A0(
        n326), .B0(n5466), .B1(n5449), .Y(n5465) );
  CLKINVX1 U7031 ( .A(n5467), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_91_N3) );
  AOI221XL U7032 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[91]), .B0(n413), .B1(N[27]), .C0(n5468), .Y(n5467) );
  OAI2B2X1 U7033 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[107]), .A0(
        n325), .B0(n5469), .B1(n5449), .Y(n5468) );
  CLKINVX1 U7034 ( .A(n5470), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_90_N3) );
  AOI221XL U7035 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[90]), .B0(n413), .B1(N[26]), .C0(n5471), .Y(n5470) );
  AO22X1 U7036 ( .A0(N[90]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[106]), .B1(n354), .Y(n5471) );
  OAI221X1 U7037 ( .A0(n5472), .A1(n369), .B0(n409), .B1(n5473), .C0(n5474), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_9_N3) );
  AOI22XL U7038 ( .A0(N[9]), .A1(n401), .B0(n350), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[25]), .Y(n5474) );
  CLKINVX1 U7039 ( .A(n5475), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_89_N3) );
  AOI221XL U7040 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[89]), .B0(n413), .B1(N[25]), .C0(n5476), .Y(n5475) );
  OAI2B2X1 U7041 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[105]), .A0(
        n326), .B0(n5477), .B1(n5449), .Y(n5476) );
  CLKINVX1 U7042 ( .A(n5478), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_88_N3) );
  AOI221XL U7043 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[88]), .B0(n413), .B1(N[24]), .C0(n5479), .Y(n5478) );
  AO22X1 U7044 ( .A0(N[88]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[104]), .B1(n354), .Y(n5479) );
  CLKINVX1 U7045 ( .A(n5480), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_87_N3) );
  AOI221XL U7046 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[87]), .B0(n413), .B1(N[23]), .C0(n5481), .Y(n5480) );
  AO22X1 U7047 ( .A0(N[87]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[79]), .B1(n354), .Y(n5481) );
  CLKINVX1 U7048 ( .A(n5482), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_86_N3) );
  AOI221XL U7049 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[86]), .B0(n413), .B1(N[22]), .C0(n5483), .Y(n5482) );
  AO22X1 U7050 ( .A0(N[86]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[78]), .B1(n354), .Y(n5483) );
  CLKINVX1 U7051 ( .A(n5484), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_85_N3) );
  AOI221XL U7052 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[85]), .B0(n413), .B1(N[21]), .C0(n5485), .Y(n5484) );
  AO22X1 U7053 ( .A0(N[85]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[77]), .B1(n354), .Y(n5485) );
  CLKINVX1 U7054 ( .A(n5486), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_84_N3) );
  AOI221XL U7055 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[84]), .B0(n413), .B1(N[20]), .C0(n5487), .Y(n5486) );
  OAI2B2X1 U7056 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[76]), .A0(n326), .B0(n5488), .B1(n5449), .Y(n5487) );
  CLKINVX1 U7057 ( .A(n5489), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_83_N3) );
  AOI221XL U7058 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[83]), .B0(n413), .B1(N[19]), .C0(n5490), .Y(n5489) );
  AO22X1 U7059 ( .A0(N[83]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[75]), .B1(n354), .Y(n5490) );
  OAI221X1 U7060 ( .A0(n364), .A1(n5491), .B0(n409), .B1(n5492), .C0(n5493), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_82_N3) );
  AOI22XL U7061 ( .A0(N[82]), .A1(n401), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[74]), .B1(n354), .Y(n5493) );
  CLKINVX1 U7062 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[82]), .Y(n5491)
         );
  CLKINVX1 U7063 ( .A(n5494), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_81_N3) );
  AOI221XL U7064 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[81]), .B0(n413), .B1(N[17]), .C0(n5495), .Y(n5494) );
  OAI2B2X1 U7065 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[73]), .A0(n325), .B0(n5473), .B1(n5449), .Y(n5495) );
  CLKINVX1 U7066 ( .A(N[81]), .Y(n5473) );
  OAI221X1 U7067 ( .A0(n365), .A1(n5454), .B0(n409), .B1(n5496), .C0(n5497), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_80_N3) );
  AOI22XL U7068 ( .A0(N[80]), .A1(n401), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[72]), .B1(n354), .Y(n5497) );
  CLKINVX1 U7069 ( .A(N[16]), .Y(n5496) );
  CLKINVX1 U7070 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[80]), .Y(n5454)
         );
  CLKINVX1 U7071 ( .A(n5498), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_8_N3) );
  AOI221XL U7072 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[8]), .A1(n5443), 
        .B0(n413), .B1(N[80]), .C0(n5499), .Y(n5498) );
  OAI2B2X1 U7073 ( .A1N(N[8]), .A0(n5449), .B0(n327), .B1(n5500), .Y(n5499) );
  CLKINVX1 U7074 ( .A(n5501), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_79_N3) );
  AOI221XL U7075 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[79]), .B0(n413), .B1(N[15]), .C0(n5502), .Y(n5501) );
  OAI2B2X1 U7076 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[95]), .A0(n326), .B0(n5503), .B1(n5449), .Y(n5502) );
  CLKINVX1 U7077 ( .A(n5504), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_78_N3) );
  AOI221XL U7078 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[78]), .B0(n413), .B1(N[14]), .C0(n5505), .Y(n5504) );
  OAI2B2X1 U7079 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[94]), .A0(n325), .B0(n5506), .B1(n5449), .Y(n5505) );
  CLKINVX1 U7080 ( .A(n5507), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_77_N3) );
  AOI221XL U7081 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[77]), .B0(n413), .B1(N[13]), .C0(n5508), .Y(n5507) );
  OAI2B2X1 U7082 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[93]), .A0(n326), .B0(n5509), .B1(n5449), .Y(n5508) );
  CLKINVX1 U7083 ( .A(n5510), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_76_N3) );
  AOI221XL U7084 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[76]), .B0(n413), .B1(N[12]), .C0(n5511), .Y(n5510) );
  OAI2B2X1 U7085 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[92]), .A0(n326), .B0(n5512), .B1(n5449), .Y(n5511) );
  CLKINVX1 U7086 ( .A(n5513), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_75_N3) );
  AOI221XL U7087 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[75]), .B0(n413), .B1(N[11]), .C0(n5514), .Y(n5513) );
  OAI2B2X1 U7088 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[91]), .A0(n325), .B0(n5515), .B1(n5449), .Y(n5514) );
  CLKINVX1 U7089 ( .A(n5516), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_74_N3) );
  AOI221XL U7090 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[74]), .B0(n413), .B1(N[10]), .C0(n5517), .Y(n5516) );
  AO22X1 U7091 ( .A0(N[74]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[90]), .B1(n354), .Y(n5517) );
  CLKINVX1 U7092 ( .A(n5518), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_73_N3) );
  AOI221XL U7093 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[73]), .B0(n413), .B1(N[9]), .C0(n5519), .Y(n5518) );
  AO22X1 U7094 ( .A0(N[73]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[89]), .B1(n354), .Y(n5519) );
  CLKINVX1 U7095 ( .A(n5520), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_72_N3) );
  AOI221XL U7096 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[72]), .B0(n413), .B1(N[8]), .C0(n5521), .Y(n5520) );
  OAI2B2X1 U7097 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[88]), .A0(n326), .B0(n5522), .B1(n5449), .Y(n5521) );
  CLKINVX1 U7098 ( .A(n5523), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_71_N3) );
  AOI221XL U7099 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[71]), .B0(n413), .B1(N[7]), .C0(n5524), .Y(n5523) );
  OAI2B2X1 U7100 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[103]), .A0(
        n326), .B0(n5525), .B1(n5449), .Y(n5524) );
  CLKINVX1 U7101 ( .A(n5526), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_70_N3) );
  AOI221XL U7102 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[70]), .B0(n413), .B1(N[6]), .C0(n5527), .Y(n5526) );
  OAI2B2X1 U7103 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[102]), .A0(
        n325), .B0(n5528), .B1(n5449), .Y(n5527) );
  OAI221X1 U7104 ( .A0(n5529), .A1(n368), .B0(n476), .B1(n410), .C0(n5530), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_7_N3) );
  AOI22XL U7105 ( .A0(N[7]), .A1(n401), .B0(n352), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[39]), .Y(n5530) );
  CLKINVX1 U7106 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[7]), .Y(n5529)
         );
  CLKINVX1 U7107 ( .A(n5531), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_69_N3) );
  AOI221XL U7108 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[69]), .B0(n413), .B1(N[5]), .C0(n5532), .Y(n5531) );
  OAI2B2X1 U7109 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[101]), .A0(
        n325), .B0(n5533), .B1(n5449), .Y(n5532) );
  CLKINVX1 U7110 ( .A(n5534), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_68_N3) );
  AOI221XL U7111 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[68]), .B0(n413), .B1(N[4]), .C0(n5535), .Y(n5534) );
  OAI2B2X1 U7112 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[100]), .A0(
        n325), .B0(n5536), .B1(n5449), .Y(n5535) );
  CLKINVX1 U7113 ( .A(n5537), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_67_N3) );
  AOI221XL U7114 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[67]), .B0(n413), .B1(N[3]), .C0(n5538), .Y(n5537) );
  OAI2B2X1 U7115 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[99]), .A0(n325), .B0(n5539), .B1(n5449), .Y(n5538) );
  CLKINVX1 U7116 ( .A(n5540), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_66_N3) );
  AOI221XL U7117 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[66]), .B0(n413), .B1(N[2]), .C0(n5541), .Y(n5540) );
  AO22X1 U7118 ( .A0(N[66]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[98]), .B1(n354), .Y(n5541) );
  CLKINVX1 U7119 ( .A(n5542), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_65_N3) );
  AOI221XL U7120 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[65]), .B0(n413), .B1(N[1]), .C0(n5543), .Y(n5542) );
  AO22X1 U7121 ( .A0(N[65]), .A1(n402), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[97]), .B1(n354), .Y(n5543) );
  CLKINVX1 U7122 ( .A(n5544), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_64_N3) );
  AOI221XL U7123 ( .A0(n5443), .A1(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[64]), .B0(n413), .B1(N[0]), .C0(n5545), .Y(n5544) );
  OAI2B2X1 U7124 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[96]), .A0(n325), .B0(n5546), .B1(n5449), .Y(n5545) );
  OAI221X1 U7125 ( .A0(n5547), .A1(n368), .B0(n484), .B1(n410), .C0(n5548), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_63_N3) );
  AOI22XL U7126 ( .A0(N[63]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[55]), .Y(n5548) );
  CLKINVX1 U7127 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[63]), .Y(n5547)
         );
  OAI221X1 U7128 ( .A0(n5549), .A1(n368), .B0(n483), .B1(n410), .C0(n5550), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_62_N3) );
  AOI22XL U7129 ( .A0(N[62]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[54]), .Y(n5550) );
  CLKINVX1 U7130 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[62]), .Y(n5549)
         );
  OAI221X1 U7131 ( .A0(n5551), .A1(n368), .B0(n482), .B1(n410), .C0(n5552), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_61_N3) );
  AOI22XL U7132 ( .A0(N[61]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[53]), .Y(n5552) );
  CLKINVX1 U7133 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[61]), .Y(n5551)
         );
  OAI221X1 U7134 ( .A0(n4855), .A1(n368), .B0(n481), .B1(n410), .C0(n5553), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_60_N3) );
  AOI22XL U7135 ( .A0(N[60]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[52]), .Y(n5553) );
  CLKINVX1 U7136 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[60]), .Y(n4855)
         );
  OAI221X1 U7137 ( .A0(n5554), .A1(n368), .B0(n475), .B1(n410), .C0(n5555), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_6_N3) );
  AOI22XL U7138 ( .A0(N[6]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[38]), .Y(n5555) );
  CLKINVX1 U7139 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[6]), .Y(n5554)
         );
  OAI221X1 U7140 ( .A0(n5556), .A1(n368), .B0(n480), .B1(n410), .C0(n5557), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_59_N3) );
  AOI22XL U7141 ( .A0(N[59]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[51]), .Y(n5557) );
  CLKINVX1 U7142 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[59]), .Y(n5556)
         );
  OAI221X1 U7143 ( .A0(n5558), .A1(n368), .B0(n479), .B1(n410), .C0(n5559), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_58_N3) );
  AOI22XL U7144 ( .A0(N[58]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[50]), .Y(n5559) );
  OAI221X1 U7145 ( .A0(n5560), .A1(n368), .B0(n478), .B1(n410), .C0(n5561), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_57_N3) );
  AOI22XL U7146 ( .A0(N[57]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[49]), .Y(n5561) );
  CLKINVX1 U7147 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[57]), .Y(n5560)
         );
  OAI221X1 U7148 ( .A0(n4895), .A1(n368), .B0(n477), .B1(n410), .C0(n5562), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_56_N3) );
  AOI22XL U7149 ( .A0(N[56]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[48]), .Y(n5562) );
  OAI221X1 U7150 ( .A0(n5563), .A1(n368), .B0(n468), .B1(n410), .C0(n5564), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_55_N3) );
  AOI22XL U7151 ( .A0(N[55]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[7]), .Y(n5564) );
  CLKINVX1 U7152 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[55]), .Y(n5563)
         );
  OAI221X1 U7153 ( .A0(n5565), .A1(n368), .B0(n467), .B1(n410), .C0(n5566), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_54_N3) );
  AOI22XL U7154 ( .A0(N[54]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[6]), .Y(n5566) );
  CLKINVX1 U7155 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[54]), .Y(n5565)
         );
  OAI221X1 U7156 ( .A0(n5567), .A1(n368), .B0(n466), .B1(n410), .C0(n5568), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_53_N3) );
  AOI22XL U7157 ( .A0(N[53]), .A1(n401), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[5]), .Y(n5568) );
  CLKINVX1 U7158 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[53]), .Y(n5567)
         );
  OAI221X1 U7159 ( .A0(n4658), .A1(n367), .B0(Inst_forkAE_LFSRInst_n51), .B1(
        n410), .C0(n5569), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_52_N3) );
  AOI22XL U7160 ( .A0(N[52]), .A1(n401), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[4]), .Y(n5569) );
  CLKINVX1 U7161 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[52]), .Y(n4658)
         );
  OAI221X1 U7162 ( .A0(n5570), .A1(n367), .B0(n1977), .B1(n410), .C0(n5571), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_51_N3) );
  AOI22XL U7163 ( .A0(N[51]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[3]), .Y(n5571) );
  CLKINVX1 U7164 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[51]), .Y(n5570)
         );
  OAI221X1 U7165 ( .A0(n5572), .A1(n367), .B0(n465), .B1(n410), .C0(n5573), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_50_N3) );
  AOI22XL U7166 ( .A0(N[50]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[2]), .Y(n5573) );
  CLKINVX1 U7167 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[50]), .Y(n5572)
         );
  OAI221X1 U7168 ( .A0(n5574), .A1(n367), .B0(n474), .B1(n410), .C0(n5575), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_5_N3) );
  AOI22XL U7169 ( .A0(N[5]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[37]), .Y(n5575) );
  CLKINVX1 U7170 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[5]), .Y(n5574)
         );
  OAI221X1 U7171 ( .A0(n5576), .A1(n367), .B0(Inst_forkAE_LFSRInst_n52), .B1(
        n409), .C0(n5577), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_49_N3) );
  AOI22XL U7172 ( .A0(N[49]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[1]), .Y(n5577) );
  CLKINVX1 U7173 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[49]), .Y(n5576)
         );
  CLKINVX1 U7174 ( .A(n5578), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_48_N3) );
  AOI221XL U7175 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[48]), .A1(n5443), .B0(Inst_forkAE_CipherInst_TK1_DEC_48_), .B1(n414), .C0(n5579), .Y(n5578) );
  OAI2B2X1 U7176 ( .A1N(N[48]), .A0(n5449), .B0(n326), .B1(n4796), .Y(n5579)
         );
  OAI221X1 U7177 ( .A0(n5580), .A1(n367), .B0(n409), .B1(n5457), .C0(n5581), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_47_N3) );
  AOI22XL U7178 ( .A0(N[47]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[63]), .Y(n5581) );
  CLKINVX1 U7179 ( .A(N[95]), .Y(n5457) );
  CLKINVX1 U7180 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[47]), .Y(n5580)
         );
  OAI221X1 U7181 ( .A0(n5582), .A1(n367), .B0(n409), .B1(n5460), .C0(n5583), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_46_N3) );
  AOI22XL U7182 ( .A0(N[46]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[62]), .Y(n5583) );
  CLKINVX1 U7183 ( .A(N[94]), .Y(n5460) );
  CLKINVX1 U7184 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[46]), .Y(n5582)
         );
  OAI221X1 U7185 ( .A0(n5584), .A1(n367), .B0(n409), .B1(n5463), .C0(n5585), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_45_N3) );
  AOI22XL U7186 ( .A0(N[45]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[61]), .Y(n5585) );
  CLKINVX1 U7187 ( .A(N[93]), .Y(n5463) );
  CLKINVX1 U7188 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[45]), .Y(n5584)
         );
  OAI221X1 U7189 ( .A0(n5586), .A1(n367), .B0(n409), .B1(n5466), .C0(n5587), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_44_N3) );
  AOI22XL U7190 ( .A0(N[44]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[60]), .Y(n5587) );
  CLKINVX1 U7191 ( .A(N[92]), .Y(n5466) );
  CLKINVX1 U7192 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[44]), .Y(n5586)
         );
  OAI221X1 U7193 ( .A0(n5588), .A1(n367), .B0(n409), .B1(n5469), .C0(n5589), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_43_N3) );
  AOI22XL U7194 ( .A0(N[43]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[59]), .Y(n5589) );
  CLKINVX1 U7195 ( .A(N[91]), .Y(n5469) );
  CLKINVX1 U7196 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[43]), .Y(n5588)
         );
  CLKINVX1 U7197 ( .A(n5590), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_42_N3) );
  AOI221XL U7198 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[42]), .A1(n5443), .B0(n413), .B1(N[90]), .C0(n5591), .Y(n5590) );
  OAI2BB2X1 U7199 ( .B0(n327), .B1(n5558), .A0N(N[42]), .A1N(n402), .Y(n5591)
         );
  CLKINVX1 U7200 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[58]), .Y(n5558)
         );
  OAI221X1 U7201 ( .A0(n5592), .A1(n369), .B0(n409), .B1(n5477), .C0(n5593), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_41_N3) );
  AOI22XL U7202 ( .A0(N[41]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[57]), .Y(n5593) );
  CLKINVX1 U7203 ( .A(N[89]), .Y(n5477) );
  CLKINVX1 U7204 ( .A(n5594), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_40_N3) );
  AOI221XL U7205 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[40]), .A1(n5443), .B0(n413), .B1(N[88]), .C0(n5595), .Y(n5594) );
  OAI2BB2X1 U7206 ( .B0(n327), .B1(n4895), .A0N(N[40]), .A1N(n402), .Y(n5595)
         );
  CLKINVX1 U7207 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[56]), .Y(n4895)
         );
  OAI221X1 U7208 ( .A0(n4756), .A1(n367), .B0(n473), .B1(n409), .C0(n5596), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_4_N3) );
  AOI22XL U7209 ( .A0(N[4]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[36]), .Y(n5596) );
  CLKINVX1 U7210 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[4]), .Y(n4756)
         );
  OAI221X1 U7211 ( .A0(n5597), .A1(n367), .B0(n409), .B1(n5525), .C0(n5598), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_39_N3) );
  AOI22XL U7212 ( .A0(N[39]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[23]), .Y(n5598) );
  CLKINVX1 U7213 ( .A(N[71]), .Y(n5525) );
  CLKINVX1 U7214 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[39]), .Y(n5597)
         );
  OAI221X1 U7215 ( .A0(n5599), .A1(n366), .B0(n408), .B1(n5528), .C0(n5600), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_38_N3) );
  AOI22XL U7216 ( .A0(N[38]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[22]), .Y(n5600) );
  CLKINVX1 U7217 ( .A(N[70]), .Y(n5528) );
  CLKINVX1 U7218 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[38]), .Y(n5599)
         );
  OAI221X1 U7219 ( .A0(n5601), .A1(n366), .B0(n408), .B1(n5533), .C0(n5602), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_37_N3) );
  AOI22XL U7220 ( .A0(N[37]), .A1(n400), .B0(n353), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[21]), .Y(n5602) );
  CLKINVX1 U7221 ( .A(N[69]), .Y(n5533) );
  CLKINVX1 U7222 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[37]), .Y(n5601)
         );
  OAI221X1 U7223 ( .A0(n5603), .A1(n366), .B0(n408), .B1(n5536), .C0(n5604), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_36_N3) );
  AOI22XL U7224 ( .A0(N[36]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[20]), .Y(n5604) );
  CLKINVX1 U7225 ( .A(N[68]), .Y(n5536) );
  CLKINVX1 U7226 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[36]), .Y(n5603)
         );
  OAI221X1 U7227 ( .A0(n5605), .A1(n366), .B0(n408), .B1(n5539), .C0(n5606), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_35_N3) );
  AOI22XL U7228 ( .A0(N[35]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[19]), .Y(n5606) );
  CLKINVX1 U7229 ( .A(N[67]), .Y(n5539) );
  CLKINVX1 U7230 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[35]), .Y(n5605)
         );
  CLKINVX1 U7231 ( .A(n5607), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_34_N3) );
  AOI221XL U7232 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[34]), .A1(n5443), .B0(n413), .B1(N[66]), .C0(n5608), .Y(n5607) );
  OAI2BB2X1 U7233 ( .B0(n327), .B1(n5609), .A0N(N[34]), .A1N(n402), .Y(n5608)
         );
  CLKINVX1 U7234 ( .A(n5610), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_33_N3) );
  AOI221XL U7235 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[33]), .A1(n5443), .B0(n413), .B1(N[65]), .C0(n5611), .Y(n5610) );
  OAI2BB2X1 U7236 ( .B0(n327), .B1(n5612), .A0N(N[33]), .A1N(n402), .Y(n5611)
         );
  OAI221X1 U7237 ( .A0(n5613), .A1(n366), .B0(n408), .B1(n5546), .C0(n5614), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_32_N3) );
  AOI22XL U7238 ( .A0(N[32]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[16]), .Y(n5614) );
  CLKINVX1 U7239 ( .A(N[64]), .Y(n5546) );
  CLKINVX1 U7240 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[32]), .Y(n5613)
         );
  OAI221X1 U7241 ( .A0(n5615), .A1(n366), .B0(n408), .B1(n5503), .C0(n5616), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_31_N3) );
  AOI22XL U7242 ( .A0(N[31]), .A1(n400), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[47]), .Y(n5616) );
  CLKINVX1 U7243 ( .A(N[79]), .Y(n5503) );
  OAI221X1 U7244 ( .A0(n5617), .A1(n366), .B0(n408), .B1(n5506), .C0(n5618), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_30_N3) );
  AOI22XL U7245 ( .A0(N[30]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[46]), .Y(n5618) );
  CLKINVX1 U7246 ( .A(N[78]), .Y(n5506) );
  OAI221X1 U7247 ( .A0(n5619), .A1(n366), .B0(n472), .B1(n409), .C0(n5620), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_3_N3) );
  AOI22XL U7248 ( .A0(N[3]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[35]), .Y(n5620) );
  CLKINVX1 U7249 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[3]), .Y(n5619)
         );
  OAI221X1 U7250 ( .A0(n5621), .A1(n366), .B0(n408), .B1(n5509), .C0(n5622), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_29_N3) );
  AOI22XL U7251 ( .A0(N[29]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[45]), .Y(n5622) );
  CLKINVX1 U7252 ( .A(N[77]), .Y(n5509) );
  OAI221X1 U7253 ( .A0(n5623), .A1(n366), .B0(n408), .B1(n5512), .C0(n5624), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_28_N3) );
  AOI22XL U7254 ( .A0(N[28]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[44]), .Y(n5624) );
  CLKINVX1 U7255 ( .A(N[76]), .Y(n5512) );
  CLKINVX1 U7256 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[28]), .Y(n5623)
         );
  OAI221X1 U7257 ( .A0(n5625), .A1(n366), .B0(n408), .B1(n5515), .C0(n5626), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_27_N3) );
  AOI22XL U7258 ( .A0(N[27]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[43]), .Y(n5626) );
  CLKINVX1 U7259 ( .A(N[75]), .Y(n5515) );
  CLKINVX1 U7260 ( .A(n5627), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_26_N3) );
  AOI221XL U7261 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[26]), .A1(n5443), .B0(n413), .B1(N[74]), .C0(n5628), .Y(n5627) );
  AO22X1 U7262 ( .A0(N[26]), .A1(n402), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[42]), .Y(n5628) );
  CLKINVX1 U7263 ( .A(n5629), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_25_N3) );
  AOI221XL U7264 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[25]), .A1(n5443), .B0(n413), .B1(N[73]), .C0(n5630), .Y(n5629) );
  OAI2BB2X1 U7265 ( .B0(n327), .B1(n5592), .A0N(N[25]), .A1N(n402), .Y(n5630)
         );
  CLKINVX1 U7266 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[41]), .Y(n5592)
         );
  OAI221X1 U7267 ( .A0(n5500), .A1(n366), .B0(n408), .B1(n5522), .C0(n5631), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_24_N3) );
  AOI22XL U7268 ( .A0(N[24]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[40]), .Y(n5631) );
  CLKINVX1 U7269 ( .A(N[72]), .Y(n5522) );
  CLKINVX1 U7270 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[24]), .Y(n5500)
         );
  CLKINVX1 U7271 ( .A(n5632), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_23_N3) );
  AOI222XL U7272 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[15]), .A1(n354), 
        .B0(n396), .B1(N[23]), .C0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[23]), .C1(n5443), .Y(n5632) );
  CLKINVX1 U7273 ( .A(n5633), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_22_N3) );
  AOI222XL U7274 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[14]), .A1(n354), 
        .B0(n395), .B1(N[22]), .C0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[22]), .C1(n5443), .Y(n5633) );
  CLKINVX1 U7275 ( .A(n5634), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_21_N3) );
  AOI222XL U7276 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[13]), .A1(n354), 
        .B0(n395), .B1(N[21]), .C0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[21]), .C1(n5443), .Y(n5634) );
  OAI211XL U7277 ( .A0(n5635), .A1(n339), .B0(n408), .C0(n5636), .Y(
        Inst_forkAE_CipherInst_KE_RS1_SFF_20_N3) );
  AOI22XL U7278 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[20]), .A1(n1989), 
        .B0(N[20]), .B1(n159), .Y(n5636) );
  OAI221X1 U7279 ( .A0(n5637), .A1(n366), .B0(n471), .B1(n409), .C0(n5638), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_2_N3) );
  AOI22XL U7280 ( .A0(N[2]), .A1(n400), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[34]), .Y(n5638) );
  CLKINVX1 U7281 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[2]), .Y(n5637)
         );
  CLKINVX1 U7282 ( .A(n5639), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_19_N3) );
  AOI222XL U7283 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[11]), .A1(n354), 
        .B0(n395), .B1(N[19]), .C0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[19]), .C1(n5443), .Y(n5639) );
  OAI222X1 U7284 ( .A0(n4311), .A1(n345), .B0(n5449), .B1(n5492), .C0(n5609), 
        .C1(n355), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_18_N3) );
  CLKINVX1 U7285 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[18]), .Y(n5609)
         );
  CLKINVX1 U7286 ( .A(N[18]), .Y(n5492) );
  OAI221X1 U7287 ( .A0(n5472), .A1(n337), .B0(n5612), .B1(n369), .C0(n5640), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_17_N3) );
  AOI32XL U7288 ( .A0(Inst_forkAE_ControlInst_fsm_state_0_), .A1(a_data), .A2(
        n414), .B0(N[17]), .B1(n399), .Y(n5640) );
  CLKINVX1 U7289 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[17]), .Y(n5612)
         );
  CLKINVX1 U7290 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[9]), .Y(n5472)
         );
  CLKINVX1 U7291 ( .A(n5641), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_16_N3) );
  AOI222XL U7292 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[8]), .A1(n354), 
        .B0(n395), .B1(N[16]), .C0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[16]), .C1(n5443), .Y(n5641) );
  CLKINVX1 U7293 ( .A(n5642), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_15_N3) );
  AOI221XL U7294 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[15]), .A1(n5443), .B0(n413), .B1(N[87]), .C0(n5643), .Y(n5642) );
  OAI2B2X1 U7295 ( .A1N(N[15]), .A0(n5449), .B0(n326), .B1(n5615), .Y(n5643)
         );
  CLKINVX1 U7296 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[31]), .Y(n5615)
         );
  CLKINVX1 U7297 ( .A(n5644), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_14_N3) );
  AOI221XL U7298 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[14]), .A1(n5443), .B0(n413), .B1(N[86]), .C0(n5645), .Y(n5644) );
  OAI2B2X1 U7299 ( .A1N(N[14]), .A0(n5449), .B0(n326), .B1(n5617), .Y(n5645)
         );
  CLKINVX1 U7300 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[30]), .Y(n5617)
         );
  CLKINVX1 U7301 ( .A(n5646), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_13_N3) );
  AOI221XL U7302 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[13]), .A1(n5443), .B0(n413), .B1(N[85]), .C0(n5647), .Y(n5646) );
  OAI2B2X1 U7303 ( .A1N(N[13]), .A0(n5449), .B0(n327), .B1(n5621), .Y(n5647)
         );
  CLKINVX1 U7304 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[29]), .Y(n5621)
         );
  CLKINVX1 U7305 ( .A(n5648), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_127_N3) );
  AOI221XL U7306 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[127]), .B0(n413), .B1(N[63]), 
        .C0(n5649), .Y(n5648) );
  OAI2BB2X1 U7307 ( .B0(n5449), .B1(n468), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[119]), .A1N(n354), .Y(n5649)
         );
  CLKINVX1 U7308 ( .A(n5650), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_126_N3) );
  AOI221XL U7309 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[126]), .B0(n413), .B1(N[62]), 
        .C0(n5651), .Y(n5650) );
  OAI2BB2X1 U7310 ( .B0(n5449), .B1(n467), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[118]), .A1N(n354), .Y(n5651)
         );
  CLKINVX1 U7311 ( .A(n5652), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_125_N3) );
  AOI221XL U7312 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[125]), .B0(n413), .B1(N[61]), 
        .C0(n5653), .Y(n5652) );
  OAI2BB2X1 U7313 ( .B0(n5449), .B1(n466), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[117]), .A1N(n354), .Y(n5653)
         );
  CLKINVX1 U7314 ( .A(n5654), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_124_N3) );
  AOI221XL U7315 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[124]), .B0(n413), .B1(N[60]), 
        .C0(n5655), .Y(n5654) );
  OAI2BB2X1 U7316 ( .B0(n5449), .B1(Inst_forkAE_LFSRInst_n51), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[116]), .A1N(n354), .Y(n5655)
         );
  CLKINVX1 U7317 ( .A(n5656), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_123_N3) );
  AOI221XL U7318 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[123]), .B0(n413), .B1(N[59]), 
        .C0(n5657), .Y(n5656) );
  OAI2B2X1 U7319 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[115]), .A0(
        n325), .B0(n5449), .B1(n1977), .Y(n5657) );
  CLKINVX1 U7320 ( .A(Inst_forkAE_CipherInst_TK1_DEC_51_), .Y(n1977) );
  CLKINVX1 U7321 ( .A(n5658), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_122_N3) );
  AOI221XL U7322 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[122]), .B0(n413), .B1(N[58]), 
        .C0(n5659), .Y(n5658) );
  OAI2BB2X1 U7323 ( .B0(n5449), .B1(n465), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[114]), .A1N(n354), .Y(n5659)
         );
  CLKINVX1 U7324 ( .A(n5660), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_121_N3) );
  AOI221XL U7325 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[121]), .B0(n413), .B1(N[57]), 
        .C0(n5661), .Y(n5660) );
  OAI2BB2X1 U7326 ( .B0(n5449), .B1(Inst_forkAE_LFSRInst_n52), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[113]), .A1N(n354), .Y(n5661)
         );
  CLKINVX1 U7327 ( .A(n5662), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_120_N3) );
  AOI221XL U7328 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[120]), .B0(n413), .B1(N[56]), 
        .C0(n5663), .Y(n5662) );
  AO22X1 U7329 ( .A0(n401), .A1(Inst_forkAE_CipherInst_TK1_DEC_48_), .B0(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[112]), .B1(n354), .Y(n5663) );
  OAI221X1 U7330 ( .A0(n5635), .A1(n365), .B0(n408), .B1(n5488), .C0(n5664), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_12_N3) );
  AOI22XL U7331 ( .A0(N[12]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[28]), .Y(n5664) );
  CLKINVX1 U7332 ( .A(N[84]), .Y(n5488) );
  CLKINVX1 U7333 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[12]), .Y(n5635)
         );
  CLKINVX1 U7334 ( .A(n5665), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_119_N3) );
  AOI221XL U7335 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[119]), .B0(n413), .B1(N[55]), 
        .C0(n5666), .Y(n5665) );
  OAI2BB2X1 U7336 ( .B0(n5449), .B1(n476), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[71]), .A1N(n354), .Y(n5666) );
  CLKINVX1 U7337 ( .A(n5667), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_118_N3) );
  AOI221XL U7338 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[118]), .B0(n413), .B1(N[54]), 
        .C0(n5668), .Y(n5667) );
  OAI2BB2X1 U7339 ( .B0(n5449), .B1(n475), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[70]), .A1N(n354), .Y(n5668) );
  CLKINVX1 U7340 ( .A(n5669), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_117_N3) );
  AOI221XL U7341 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[117]), .B0(n413), .B1(N[53]), 
        .C0(n5670), .Y(n5669) );
  OAI2BB2X1 U7342 ( .B0(n5449), .B1(n474), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[69]), .A1N(n354), .Y(n5670) );
  CLKINVX1 U7343 ( .A(n5671), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_116_N3) );
  AOI221XL U7344 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[116]), .B0(n413), .B1(N[52]), 
        .C0(n5672), .Y(n5671) );
  OAI2BB2X1 U7345 ( .B0(n5449), .B1(n473), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[68]), .A1N(n354), .Y(n5672) );
  CLKINVX1 U7346 ( .A(n5673), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_115_N3) );
  AOI221XL U7347 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[115]), .B0(n414), .B1(N[51]), 
        .C0(n5674), .Y(n5673) );
  OAI2BB2X1 U7348 ( .B0(n5449), .B1(n472), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[67]), .A1N(n354), .Y(n5674) );
  CLKINVX1 U7349 ( .A(n5675), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_114_N3) );
  AOI221XL U7350 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[114]), .B0(n414), .B1(N[50]), 
        .C0(n5676), .Y(n5675) );
  OAI2BB2X1 U7351 ( .B0(n5449), .B1(n471), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[66]), .A1N(n354), .Y(n5676) );
  CLKINVX1 U7352 ( .A(n5677), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_113_N3) );
  AOI221XL U7353 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[113]), .B0(n414), .B1(N[49]), 
        .C0(n5678), .Y(n5677) );
  OAI2BB2X1 U7354 ( .B0(n5449), .B1(n470), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[65]), .A1N(n354), .Y(n5678) );
  CLKINVX1 U7355 ( .A(n5679), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_112_N3) );
  AOI221XL U7356 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[112]), .B0(n414), .B1(N[48]), 
        .C0(n5680), .Y(n5679) );
  OAI2BB2X1 U7357 ( .B0(n5449), .B1(n469), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[64]), .A1N(n354), .Y(n5680) );
  CLKINVX1 U7358 ( .A(n5681), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_111_N3) );
  AOI221XL U7359 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[111]), .B0(n414), .B1(N[47]), 
        .C0(n5682), .Y(n5681) );
  OAI2B2X1 U7360 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[127]), .A0(
        n325), .B0(n5449), .B1(n484), .Y(n5682) );
  CLKINVX1 U7361 ( .A(n5683), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_110_N3) );
  AOI221XL U7362 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[110]), .B0(n414), .B1(N[46]), 
        .C0(n5684), .Y(n5683) );
  OAI2BB2X1 U7363 ( .B0(n5449), .B1(n483), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[126]), .A1N(n354), .Y(n5684)
         );
  CLKINVX1 U7364 ( .A(n5685), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_11_N3) );
  AOI221XL U7365 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[11]), .A1(n5443), .B0(n414), .B1(N[83]), .C0(n5686), .Y(n5685) );
  OAI2B2X1 U7366 ( .A1N(N[11]), .A0(n5449), .B0(n326), .B1(n5625), .Y(n5686)
         );
  CLKINVX1 U7367 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[27]), .Y(n5625)
         );
  CLKINVX1 U7368 ( .A(n5687), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_109_N3) );
  AOI221XL U7369 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[109]), .B0(n414), .B1(N[45]), 
        .C0(n5688), .Y(n5687) );
  OAI2BB2X1 U7370 ( .B0(n5449), .B1(n482), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[125]), .A1N(n354), .Y(n5688)
         );
  CLKINVX1 U7371 ( .A(n5689), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_108_N3) );
  AOI221XL U7372 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[108]), .B0(n414), .B1(N[44]), 
        .C0(n5690), .Y(n5689) );
  OAI2BB2X1 U7373 ( .B0(n5449), .B1(n481), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[124]), .A1N(n354), .Y(n5690)
         );
  CLKINVX1 U7374 ( .A(n5691), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_107_N3) );
  AOI221XL U7375 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[107]), .B0(n414), .B1(N[43]), 
        .C0(n5692), .Y(n5691) );
  OAI2BB2X1 U7376 ( .B0(n5449), .B1(n480), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[123]), .A1N(n354), .Y(n5692)
         );
  CLKINVX1 U7377 ( .A(n5693), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_106_N3) );
  AOI221XL U7378 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[106]), .B0(n414), .B1(N[42]), 
        .C0(n5694), .Y(n5693) );
  OAI2BB2X1 U7379 ( .B0(n5449), .B1(n479), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[122]), .A1N(n354), .Y(n5694)
         );
  CLKINVX1 U7380 ( .A(n5695), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_105_N3) );
  AOI221XL U7381 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[105]), .B0(n414), .B1(N[41]), 
        .C0(n5696), .Y(n5695) );
  OAI2BB2X1 U7382 ( .B0(n5449), .B1(n478), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[121]), .A1N(n354), .Y(n5696)
         );
  CLKINVX1 U7383 ( .A(n5697), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_104_N3) );
  AOI221XL U7384 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[104]), .B0(n414), .B1(N[40]), 
        .C0(n5698), .Y(n5697) );
  OAI2BB2X1 U7385 ( .B0(n5449), .B1(n477), .A0N(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[120]), .A1N(n354), .Y(n5698)
         );
  CLKINVX1 U7386 ( .A(n5699), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_103_N3) );
  AOI222XL U7387 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[103]), .B0(n349), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[87]), .C0(n414), .C1(N[39]), 
        .Y(n5699) );
  CLKINVX1 U7388 ( .A(n5700), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_102_N3) );
  AOI222XL U7389 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[102]), .B0(n346), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[86]), .C0(n414), .C1(N[38]), 
        .Y(n5700) );
  CLKINVX1 U7390 ( .A(n5701), .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_101_N3) );
  AOI222XL U7391 ( .A0(n5443), .A1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[101]), .B0(n348), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[85]), .C0(n414), .C1(N[37]), 
        .Y(n5701) );
  OAI2B11X1 U7392 ( .A1N(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[100]), .A0(
        n355), .B0(n5449), .C0(n5702), .Y(
        Inst_forkAE_CipherInst_KE_RS1_SFF_100_N3) );
  AOI22XL U7393 ( .A0(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[84]), .A1(n2244), 
        .B0(N[36]), .B1(n159), .Y(n5702) );
  OAI221X1 U7394 ( .A0(n4311), .A1(n367), .B0(n408), .B1(n5703), .C0(n5704), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_10_N3) );
  AOI22XL U7395 ( .A0(N[10]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[26]), .Y(n5704) );
  CLKINVX1 U7396 ( .A(N[82]), .Y(n5703) );
  CLKINVX1 U7397 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[10]), .Y(n4311)
         );
  OAI221X1 U7398 ( .A0(n5705), .A1(n365), .B0(n470), .B1(n409), .C0(n5706), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_1_N3) );
  AOI22XL U7399 ( .A0(N[1]), .A1(n399), .B0(n354), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[33]), .Y(n5706) );
  CLKINVX1 U7400 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[1]), .Y(n5705)
         );
  OAI221X1 U7401 ( .A0(n4796), .A1(n365), .B0(n469), .B1(n409), .C0(n5707), 
        .Y(Inst_forkAE_CipherInst_KE_RS1_SFF_0_N3) );
  AOI22XL U7402 ( .A0(N[0]), .A1(n399), .B0(n351), .B1(
        Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[32]), .Y(n5707) );
  CLKINVX1 U7403 ( .A(n5449), .Y(n5192) );
  CLKNAND2X2 U7404 ( .A(n2244), .B(n145), .Y(n5449) );
  CLKINVX1 U7405 ( .A(n5443), .Y(n4963) );
  CLKINVX1 U7406 ( .A(Inst_forkAE_CipherInst_KE_KEY_PERM1_Inv[0]), .Y(n4796)
         );
  NOR2BX1 U7407 ( .AN(clk), .B(n462), .Y(Inst_forkAE_CipherInst_KE_CLK_K) );
  CLKNAND2X2 U7408 ( .A(n5708), .B(n408), .Y(Inst_forkAE_CipherInst_CL_n44) );
  MXI2X1 U7409 ( .A(n5709), .B(Inst_forkAE_CipherInst_CL_STATE_0_), .S0(
        Inst_forkAE_CipherInst_CL_n34), .Y(n5708) );
  NOR2X1 U7410 ( .A(n1996), .B(n145), .Y(n5709) );
  MXI2X1 U7411 ( .A(n5710), .B(n464), .S0(n1989), .Y(n1996) );
  XOR2X1 U7412 ( .A(n4), .B(Inst_forkAE_CipherInst_CL_n23), .Y(n5710) );
  CLKNAND2X2 U7413 ( .A(n5711), .B(n408), .Y(Inst_forkAE_CipherInst_CL_n43) );
  MXI2X1 U7414 ( .A(n5712), .B(n461), .S0(Inst_forkAE_CipherInst_CL_n34), .Y(
        n5711) );
  NOR2X1 U7415 ( .A(n4670), .B(n145), .Y(n5712) );
  CLKINVX1 U7416 ( .A(Inst_forkAE_ControlInst_fsm_state_1_), .Y(n1985) );
  CLKINVX1 U7417 ( .A(n1994), .Y(n4670) );
  MXI2X1 U7418 ( .A(Inst_forkAE_CipherInst_CL_n27), .B(
        Inst_forkAE_CipherInst_CL_n23), .S0(n1989), .Y(n1994) );
  CLKINVX1 U7419 ( .A(n2288), .Y(n2254) );
  CLKINVX1 U7420 ( .A(n4584), .Y(n3977) );
  CLKNAND2X2 U7421 ( .A(Block_Size[1]), .B(n4495), .Y(n4584) );
  CLKINVX1 U7422 ( .A(n4322), .Y(n4495) );
  CLKNAND2X2 U7423 ( .A(Block_Size[3]), .B(Block_Size[2]), .Y(n4322) );
  MXI2X1 U7424 ( .A(n5713), .B(n5714), .S0(
        Inst_forkAE_CipherInst_CL_COUNTER_2_), .Y(
        Inst_forkAE_CipherInst_CL_N15) );
  AOI21X1 U7425 ( .A0(n463), .A1(Inst_forkAE_CipherInst_CL_n34), .B0(
        Inst_forkAE_CipherInst_CL_N13), .Y(n5714) );
  NAND3XL U7426 ( .A(Inst_forkAE_CipherInst_CL_n34), .B(n2), .C(
        Inst_forkAE_CipherInst_CL_COUNTER_0_), .Y(n5713) );
  CLKINVX1 U7427 ( .A(Inst_forkAE_CipherInst_KE_N2), .Y(
        Inst_forkAE_CipherInst_CL_n34) );
  NOR2X1 U7428 ( .A(Inst_forkAE_CipherInst_KE_N2), .B(
        Inst_forkAE_CipherInst_CL_COUNTER_0_), .Y(
        Inst_forkAE_CipherInst_CL_N13) );
  CLKNAND2X2 U7429 ( .A(Inst_forkAE_ControlInst_fsm_state_1_), .B(n1993), .Y(
        Inst_forkAE_CipherInst_KE_N2) );
  CLKINVX1 U7430 ( .A(Inst_forkAE_CipherInst_LAST), .Y(n1993) );
  NOR3BX1 U7431 ( .AN(Inst_forkAE_CipherInst_CL_COUNTER_2_), .B(
        Inst_forkAE_CipherInst_CL_COUNTER_0_), .C(n2), .Y(
        Inst_forkAE_CipherInst_LAST) );
endmodule


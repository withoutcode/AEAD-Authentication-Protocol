
module forkAE_imp ( clk, rst, en_c, ld_rec, IDt, IDst, key, DtSel, rand_in, 
        MuxSel2, GO, ENC_DEC_MODE, DONE, PLAINTEXT, C1, C0 );
  input [63:0] IDt;
  input [63:0] IDst;
  input [127:0] key;
  input [63:0] rand_in;
  input [63:0] PLAINTEXT;
  output [63:0] C1;
  output [63:0] C0;
  input clk, rst, en_c, ld_rec, DtSel, MuxSel2, GO, ENC_DEC_MODE;
  output DONE;
  wire   Inst_forkAE_CURRENT_KEY_35_, Inst_forkAE_CURRENT_KEY_39_,
         Inst_forkAE_CURRENT_KEY_43_, Inst_forkAE_CURRENT_KEY_47_,
         Inst_forkAE_CURRENT_KEY_51_, Inst_forkAE_CURRENT_KEY_55_,
         Inst_forkAE_CURRENT_KEY_59_, Inst_forkAE_CURRENT_KEY_63_,
         Inst_forkAE_CURRENT_KEY_96_, Inst_forkAE_CURRENT_KEY_100_,
         Inst_forkAE_CURRENT_KEY_104_, Inst_forkAE_CURRENT_KEY_108_,
         Inst_forkAE_CURRENT_KEY_112_, Inst_forkAE_CURRENT_KEY_116_,
         Inst_forkAE_CURRENT_KEY_120_, Inst_forkAE_CURRENT_KEY_124_,
         Inst_forkAE_CONST_ENC_1_, Inst_forkAE_CONST_ENC_2_,
         Inst_forkAE_CONST_ENC_5_, Inst_forkAE_CONST_DEC_6_, Inst_lfsr_n195,
         Inst_lfsr_n194, Inst_lfsr_n193, Inst_lfsr_n192, Inst_lfsr_n191,
         Inst_lfsr_n190, Inst_lfsr_n189, Inst_lfsr_n188, Inst_lfsr_n187,
         Inst_lfsr_n186, Inst_lfsr_n185, Inst_lfsr_n184, Inst_lfsr_n183,
         Inst_lfsr_n182, Inst_lfsr_n181, Inst_lfsr_n180, Inst_lfsr_n179,
         Inst_lfsr_n178, Inst_lfsr_n177, Inst_lfsr_n176, Inst_lfsr_n175,
         Inst_lfsr_n174, Inst_lfsr_n173, Inst_lfsr_n172, Inst_lfsr_n171,
         Inst_lfsr_n170, Inst_lfsr_n169, Inst_lfsr_n168, Inst_lfsr_n167,
         Inst_lfsr_n166, Inst_lfsr_n165, Inst_lfsr_n164, Inst_lfsr_n163,
         Inst_lfsr_n162, Inst_lfsr_n161, Inst_lfsr_n160, Inst_lfsr_n159,
         Inst_lfsr_n158, Inst_lfsr_n157, Inst_lfsr_n156, Inst_lfsr_n155,
         Inst_lfsr_n154, Inst_lfsr_n153, Inst_lfsr_n152, Inst_lfsr_n151,
         Inst_lfsr_n150, Inst_lfsr_n149, Inst_lfsr_n148, Inst_lfsr_n147,
         Inst_lfsr_n146, Inst_lfsr_n145, Inst_lfsr_n144, Inst_lfsr_n143,
         Inst_lfsr_n142, Inst_lfsr_n141, Inst_lfsr_n140, Inst_lfsr_n139,
         Inst_lfsr_n138, Inst_lfsr_n137, Inst_lfsr_n136, Inst_lfsr_n135,
         Inst_lfsr_n134, Inst_lfsr_n133, Inst_lfsr_n132, Inst_lfsr_N66,
         Inst_lfsr_N65, Inst_lfsr_N64, Inst_lfsr_N63, Inst_lfsr_N62,
         Inst_lfsr_N61, Inst_lfsr_N60, Inst_lfsr_N59, Inst_lfsr_N58,
         Inst_lfsr_N57, Inst_lfsr_N56, Inst_lfsr_N55, Inst_lfsr_N54,
         Inst_lfsr_N53, Inst_lfsr_N52, Inst_lfsr_N51, Inst_lfsr_N50,
         Inst_lfsr_N49, Inst_lfsr_N48, Inst_lfsr_N47, Inst_lfsr_N46,
         Inst_lfsr_N45, Inst_lfsr_N44, Inst_lfsr_N43, Inst_lfsr_N42,
         Inst_lfsr_N41, Inst_lfsr_N40, Inst_lfsr_N39, Inst_lfsr_N38,
         Inst_lfsr_N37, Inst_lfsr_N36, Inst_lfsr_N35, Inst_lfsr_N34,
         Inst_lfsr_N33, Inst_lfsr_N32, Inst_lfsr_N31, Inst_lfsr_N30,
         Inst_lfsr_N29, Inst_lfsr_N28, Inst_lfsr_N27, Inst_lfsr_N26,
         Inst_lfsr_N25, Inst_lfsr_N24, Inst_lfsr_N23, Inst_lfsr_N22,
         Inst_lfsr_N21, Inst_lfsr_N20, Inst_lfsr_N19, Inst_lfsr_N18,
         Inst_lfsr_N17, Inst_lfsr_N16, Inst_lfsr_N15, Inst_lfsr_N14,
         Inst_lfsr_N13, Inst_lfsr_N12, Inst_lfsr_N11, Inst_lfsr_N10,
         Inst_lfsr_N9, Inst_lfsr_N8, Inst_lfsr_N7, Inst_lfsr_N6, Inst_lfsr_N5,
         Inst_RegIDt_n130, Inst_RegIDt_n127, Inst_RegIDt_n125,
         Inst_RegIDt_n123, Inst_RegIDt_n121, Inst_RegIDt_n119,
         Inst_RegIDt_n117, Inst_RegIDt_n115, Inst_RegIDt_n113,
         Inst_RegIDt_n111, Inst_RegIDt_n109, Inst_RegIDt_n107,
         Inst_RegIDt_n105, Inst_RegIDt_n103, Inst_RegIDt_n101, Inst_RegIDt_n99,
         Inst_RegIDt_n97, Inst_RegIDt_n95, Inst_RegIDt_n93, Inst_RegIDt_n91,
         Inst_RegIDt_n89, Inst_RegIDt_n87, Inst_RegIDt_n85, Inst_RegIDt_n83,
         Inst_RegIDt_n81, Inst_RegIDt_n79, Inst_RegIDt_n77, Inst_RegIDt_n75,
         Inst_RegIDt_n73, Inst_RegIDt_n71, Inst_RegIDt_n69, Inst_RegIDt_n67,
         Inst_RegIDt_n65, Inst_RegIDt_n63, Inst_RegIDt_n61, Inst_RegIDt_n59,
         Inst_RegIDt_n57, Inst_RegIDt_n55, Inst_RegIDt_n53, Inst_RegIDt_n51,
         Inst_RegIDt_n49, Inst_RegIDt_n47, Inst_RegIDt_n45, Inst_RegIDt_n43,
         Inst_RegIDt_n41, Inst_RegIDt_n39, Inst_RegIDt_n37, Inst_RegIDt_n35,
         Inst_RegIDt_n33, Inst_RegIDt_n31, Inst_RegIDt_n29, Inst_RegIDt_n27,
         Inst_RegIDt_n25, Inst_RegIDt_n23, Inst_RegIDt_n21, Inst_RegIDt_n19,
         Inst_RegIDt_n17, Inst_RegIDt_n15, Inst_RegIDt_n13, Inst_RegIDt_n11,
         Inst_RegIDt_n9, Inst_RegIDt_n7, Inst_RegIDt_n5, Inst_RegIDt_n3,
         Inst_forkAE_FSM_X_N43, Inst_forkAE_FSM_X_N42, Inst_forkAE_FSM_X_N41,
         Inst_forkAE_FSM_X_state_0_, Inst_forkAE_FSM_X_state_1_,
         Inst_forkAE_FSM_X_state_2_, Inst_forkAE_REG_INTERNAL_STATE_N65,
         Inst_forkAE_REG_INTERNAL_STATE_N64,
         Inst_forkAE_REG_INTERNAL_STATE_N63,
         Inst_forkAE_REG_INTERNAL_STATE_N62,
         Inst_forkAE_REG_INTERNAL_STATE_N61,
         Inst_forkAE_REG_INTERNAL_STATE_N60,
         Inst_forkAE_REG_INTERNAL_STATE_N59,
         Inst_forkAE_REG_INTERNAL_STATE_N58,
         Inst_forkAE_REG_INTERNAL_STATE_N57,
         Inst_forkAE_REG_INTERNAL_STATE_N56,
         Inst_forkAE_REG_INTERNAL_STATE_N55,
         Inst_forkAE_REG_INTERNAL_STATE_N54,
         Inst_forkAE_REG_INTERNAL_STATE_N53,
         Inst_forkAE_REG_INTERNAL_STATE_N52,
         Inst_forkAE_REG_INTERNAL_STATE_N51,
         Inst_forkAE_REG_INTERNAL_STATE_N50,
         Inst_forkAE_REG_INTERNAL_STATE_N49,
         Inst_forkAE_REG_INTERNAL_STATE_N48,
         Inst_forkAE_REG_INTERNAL_STATE_N47,
         Inst_forkAE_REG_INTERNAL_STATE_N46,
         Inst_forkAE_REG_INTERNAL_STATE_N45,
         Inst_forkAE_REG_INTERNAL_STATE_N44,
         Inst_forkAE_REG_INTERNAL_STATE_N43,
         Inst_forkAE_REG_INTERNAL_STATE_N42,
         Inst_forkAE_REG_INTERNAL_STATE_N41,
         Inst_forkAE_REG_INTERNAL_STATE_N40,
         Inst_forkAE_REG_INTERNAL_STATE_N39,
         Inst_forkAE_REG_INTERNAL_STATE_N38,
         Inst_forkAE_REG_INTERNAL_STATE_N37,
         Inst_forkAE_REG_INTERNAL_STATE_N36,
         Inst_forkAE_REG_INTERNAL_STATE_N35,
         Inst_forkAE_REG_INTERNAL_STATE_N34,
         Inst_forkAE_REG_INTERNAL_STATE_N33,
         Inst_forkAE_REG_INTERNAL_STATE_N32,
         Inst_forkAE_REG_INTERNAL_STATE_N31,
         Inst_forkAE_REG_INTERNAL_STATE_N30,
         Inst_forkAE_REG_INTERNAL_STATE_N29,
         Inst_forkAE_REG_INTERNAL_STATE_N28,
         Inst_forkAE_REG_INTERNAL_STATE_N27,
         Inst_forkAE_REG_INTERNAL_STATE_N26,
         Inst_forkAE_REG_INTERNAL_STATE_N25,
         Inst_forkAE_REG_INTERNAL_STATE_N24,
         Inst_forkAE_REG_INTERNAL_STATE_N23,
         Inst_forkAE_REG_INTERNAL_STATE_N22,
         Inst_forkAE_REG_INTERNAL_STATE_N21,
         Inst_forkAE_REG_INTERNAL_STATE_N20,
         Inst_forkAE_REG_INTERNAL_STATE_N19,
         Inst_forkAE_REG_INTERNAL_STATE_N18,
         Inst_forkAE_REG_INTERNAL_STATE_N17,
         Inst_forkAE_REG_INTERNAL_STATE_N16,
         Inst_forkAE_REG_INTERNAL_STATE_N15,
         Inst_forkAE_REG_INTERNAL_STATE_N14,
         Inst_forkAE_REG_INTERNAL_STATE_N13,
         Inst_forkAE_REG_INTERNAL_STATE_N12,
         Inst_forkAE_REG_INTERNAL_STATE_N11,
         Inst_forkAE_REG_INTERNAL_STATE_N10, Inst_forkAE_REG_INTERNAL_STATE_N9,
         Inst_forkAE_REG_INTERNAL_STATE_N8, Inst_forkAE_REG_INTERNAL_STATE_N7,
         Inst_forkAE_REG_INTERNAL_STATE_N6, Inst_forkAE_REG_INTERNAL_STATE_N5,
         Inst_forkAE_REG_INTERNAL_STATE_N4, Inst_forkAE_REG_INTERNAL_STATE_N3,
         Inst_forkAE_REG_INTERNAL_STATE_N2, Inst_forkAE_ConstGen_N30,
         Inst_forkAE_ConstGen_N28, Inst_forkAE_ConstGen_N25,
         Inst_forkAE_ConstGen_N24, Inst_forkAE_REG_TK2_0_N65,
         Inst_forkAE_REG_TK2_0_N64, Inst_forkAE_REG_TK2_0_N63,
         Inst_forkAE_REG_TK2_0_N62, Inst_forkAE_REG_TK2_0_N61,
         Inst_forkAE_REG_TK2_0_N60, Inst_forkAE_REG_TK2_0_N59,
         Inst_forkAE_REG_TK2_0_N58, Inst_forkAE_REG_TK2_0_N57,
         Inst_forkAE_REG_TK2_0_N56, Inst_forkAE_REG_TK2_0_N55,
         Inst_forkAE_REG_TK2_0_N54, Inst_forkAE_REG_TK2_0_N53,
         Inst_forkAE_REG_TK2_0_N52, Inst_forkAE_REG_TK2_0_N51,
         Inst_forkAE_REG_TK2_0_N50, Inst_forkAE_REG_TK2_0_N49,
         Inst_forkAE_REG_TK2_0_N48, Inst_forkAE_REG_TK2_0_N47,
         Inst_forkAE_REG_TK2_0_N46, Inst_forkAE_REG_TK2_0_N45,
         Inst_forkAE_REG_TK2_0_N44, Inst_forkAE_REG_TK2_0_N43,
         Inst_forkAE_REG_TK2_0_N42, Inst_forkAE_REG_TK2_0_N41,
         Inst_forkAE_REG_TK2_0_N40, Inst_forkAE_REG_TK2_0_N39,
         Inst_forkAE_REG_TK2_0_N38, Inst_forkAE_REG_TK2_0_N37,
         Inst_forkAE_REG_TK2_0_N36, Inst_forkAE_REG_TK2_0_N35,
         Inst_forkAE_REG_TK2_0_N34, Inst_forkAE_REG_TK2_0_N33,
         Inst_forkAE_REG_TK2_0_N32, Inst_forkAE_REG_TK2_0_N31,
         Inst_forkAE_REG_TK2_0_N30, Inst_forkAE_REG_TK2_0_N29,
         Inst_forkAE_REG_TK2_0_N28, Inst_forkAE_REG_TK2_0_N27,
         Inst_forkAE_REG_TK2_0_N26, Inst_forkAE_REG_TK2_0_N25,
         Inst_forkAE_REG_TK2_0_N24, Inst_forkAE_REG_TK2_0_N23,
         Inst_forkAE_REG_TK2_0_N22, Inst_forkAE_REG_TK2_0_N21,
         Inst_forkAE_REG_TK2_0_N20, Inst_forkAE_REG_TK2_0_N19,
         Inst_forkAE_REG_TK2_0_N18, Inst_forkAE_REG_TK2_0_N17,
         Inst_forkAE_REG_TK2_0_N16, Inst_forkAE_REG_TK2_0_N15,
         Inst_forkAE_REG_TK2_0_N14, Inst_forkAE_REG_TK2_0_N13,
         Inst_forkAE_REG_TK2_0_N12, Inst_forkAE_REG_TK2_0_N11,
         Inst_forkAE_REG_TK2_0_N10, Inst_forkAE_REG_TK2_0_N9,
         Inst_forkAE_REG_TK2_0_N8, Inst_forkAE_REG_TK2_0_N7,
         Inst_forkAE_REG_TK2_0_N6, Inst_forkAE_REG_TK2_0_N5,
         Inst_forkAE_REG_TK2_0_N4, Inst_forkAE_REG_TK2_0_N3,
         Inst_forkAE_REG_TK2_0_N2, Inst_forkAE_REG_TK2_N65,
         Inst_forkAE_REG_TK2_N64, Inst_forkAE_REG_TK2_N63,
         Inst_forkAE_REG_TK2_N62, Inst_forkAE_REG_TK2_N61,
         Inst_forkAE_REG_TK2_N60, Inst_forkAE_REG_TK2_N59,
         Inst_forkAE_REG_TK2_N58, Inst_forkAE_REG_TK2_N57,
         Inst_forkAE_REG_TK2_N56, Inst_forkAE_REG_TK2_N55,
         Inst_forkAE_REG_TK2_N54, Inst_forkAE_REG_TK2_N53,
         Inst_forkAE_REG_TK2_N52, Inst_forkAE_REG_TK2_N51,
         Inst_forkAE_REG_TK2_N50, Inst_forkAE_REG_TK2_N49,
         Inst_forkAE_REG_TK2_N48, Inst_forkAE_REG_TK2_N47,
         Inst_forkAE_REG_TK2_N46, Inst_forkAE_REG_TK2_N45,
         Inst_forkAE_REG_TK2_N44, Inst_forkAE_REG_TK2_N43,
         Inst_forkAE_REG_TK2_N42, Inst_forkAE_REG_TK2_N41,
         Inst_forkAE_REG_TK2_N40, Inst_forkAE_REG_TK2_N39,
         Inst_forkAE_REG_TK2_N38, Inst_forkAE_REG_TK2_N37,
         Inst_forkAE_REG_TK2_N36, Inst_forkAE_REG_TK2_N35,
         Inst_forkAE_REG_TK2_N34, Inst_forkAE_REG_TK2_N33,
         Inst_forkAE_REG_TK2_N32, Inst_forkAE_REG_TK2_N31,
         Inst_forkAE_REG_TK2_N30, Inst_forkAE_REG_TK2_N29,
         Inst_forkAE_REG_TK2_N28, Inst_forkAE_REG_TK2_N27,
         Inst_forkAE_REG_TK2_N26, Inst_forkAE_REG_TK2_N25,
         Inst_forkAE_REG_TK2_N24, Inst_forkAE_REG_TK2_N23,
         Inst_forkAE_REG_TK2_N22, Inst_forkAE_REG_TK2_N21,
         Inst_forkAE_REG_TK2_N20, Inst_forkAE_REG_TK2_N19,
         Inst_forkAE_REG_TK2_N18, Inst_forkAE_REG_TK2_N17,
         Inst_forkAE_REG_TK2_N16, Inst_forkAE_REG_TK2_N15,
         Inst_forkAE_REG_TK2_N14, Inst_forkAE_REG_TK2_N13,
         Inst_forkAE_REG_TK2_N12, Inst_forkAE_REG_TK2_N11,
         Inst_forkAE_REG_TK2_N10, Inst_forkAE_REG_TK2_N9,
         Inst_forkAE_REG_TK2_N8, Inst_forkAE_REG_TK2_N7,
         Inst_forkAE_REG_TK2_N6, Inst_forkAE_REG_TK2_N5,
         Inst_forkAE_REG_TK2_N4, Inst_forkAE_REG_TK2_N3,
         Inst_forkAE_REG_TK2_N2, Inst_forkAE_L_N65, Inst_forkAE_L_N64,
         Inst_forkAE_L_N63, Inst_forkAE_L_N62, Inst_forkAE_L_N61,
         Inst_forkAE_L_N60, Inst_forkAE_L_N59, Inst_forkAE_L_N58,
         Inst_forkAE_L_N57, Inst_forkAE_L_N56, Inst_forkAE_L_N55,
         Inst_forkAE_L_N54, Inst_forkAE_L_N53, Inst_forkAE_L_N52,
         Inst_forkAE_L_N51, Inst_forkAE_L_N50, Inst_forkAE_L_N49,
         Inst_forkAE_L_N48, Inst_forkAE_L_N47, Inst_forkAE_L_N46,
         Inst_forkAE_L_N45, Inst_forkAE_L_N44, Inst_forkAE_L_N43,
         Inst_forkAE_L_N42, Inst_forkAE_L_N41, Inst_forkAE_L_N40,
         Inst_forkAE_L_N39, Inst_forkAE_L_N38, Inst_forkAE_L_N37,
         Inst_forkAE_L_N36, Inst_forkAE_L_N35, Inst_forkAE_L_N34,
         Inst_forkAE_L_N33, Inst_forkAE_L_N32, Inst_forkAE_L_N31,
         Inst_forkAE_L_N30, Inst_forkAE_L_N29, Inst_forkAE_L_N28,
         Inst_forkAE_L_N27, Inst_forkAE_L_N26, Inst_forkAE_L_N25,
         Inst_forkAE_L_N24, Inst_forkAE_L_N23, Inst_forkAE_L_N22,
         Inst_forkAE_L_N21, Inst_forkAE_L_N20, Inst_forkAE_L_N19,
         Inst_forkAE_L_N18, Inst_forkAE_L_N17, Inst_forkAE_L_N16,
         Inst_forkAE_L_N15, Inst_forkAE_L_N14, Inst_forkAE_L_N13,
         Inst_forkAE_L_N12, Inst_forkAE_L_N11, Inst_forkAE_L_N10,
         Inst_forkAE_L_N9, Inst_forkAE_L_N8, Inst_forkAE_L_N7,
         Inst_forkAE_L_N6, Inst_forkAE_L_N5, Inst_forkAE_L_N4,
         Inst_forkAE_L_N3, Inst_forkAE_L_N2, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2622, n2624, n2626, n2628, n2630, n2632,
         n2634, n2636, n2638, n2640, n2642, n2644, n2646, n2648, n2650, n2652,
         n2654, n2656, n2658, n2660, n2662, n2664, n2666, n2668, n2670, n2672,
         n2674, n2676, n2678, n2680, n2682, n2684, n2686, n2688, n2690, n2692,
         n2694, n2696, n2698, n2700, n2702, n2704, n2706, n2708, n2710, n2712,
         n2714, n2716, n2718, n2720, n2722, n2724, n2726, n2728, n2730, n2732,
         n2734, n2736, n2738, n2740, n2742, n2744, n2746, n2748;
  wire   [63:0] randd;
  wire   [63:0] IDtReg;
  wire   [63:0] IDstReg;
  wire   [191:1] Inst_forkAE_KEY_INVERSE;
  wire   [63:2] Inst_lfsr_add_3205_carry;

  SDFFTRXL Inst_forkAE_ConstGen_STATE_reg_5_ ( .RN(Inst_forkAE_FSM_X_state_0_), 
        .D(n2106), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n131), .QN(n181) );
  SDFFTRXL Inst_forkAE_ConstGen_STATE_reg_3_ ( .RN(Inst_forkAE_FSM_X_state_0_), 
        .D(n2107), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n133), .QN(n180) );
  SDFFTRXL Inst_forkAE_ConstGen_STATE_reg_2_ ( .RN(Inst_forkAE_FSM_X_state_0_), 
        .D(n2108), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n132), .QN(n179) );
  SDFFSQXL Inst_forkAE_L_Q_reg_4_ ( .D(Inst_forkAE_L_N6), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[4]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_12_ ( .D(Inst_forkAE_L_N14), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[12]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_40_ ( .D(Inst_forkAE_L_N42), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[40]) );
  SDFFRQX2 Inst_REgIDst_do_reg_0_ ( .D(n2622), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[0]) );
  SDFFRQX2 Inst_REgIDst_do_reg_1_ ( .D(n2624), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[1]) );
  SDFFRQX2 Inst_REgIDst_do_reg_2_ ( .D(n2626), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[2]) );
  SDFFRQX2 Inst_REgIDst_do_reg_3_ ( .D(n2628), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[3]) );
  SDFFRQX2 Inst_REgIDst_do_reg_4_ ( .D(n2630), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[4]) );
  SDFFRQX2 Inst_REgIDst_do_reg_5_ ( .D(n2632), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[5]) );
  SDFFRQX2 Inst_REgIDst_do_reg_6_ ( .D(n2634), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[6]) );
  SDFFRQX2 Inst_REgIDst_do_reg_7_ ( .D(n2636), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n169), .Q(IDstReg[7]) );
  SDFFRQX2 Inst_REgIDst_do_reg_8_ ( .D(n2638), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[8]) );
  SDFFRQX2 Inst_REgIDst_do_reg_9_ ( .D(n2640), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[9]) );
  SDFFRQX2 Inst_REgIDst_do_reg_10_ ( .D(n2642), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[10]) );
  SDFFRQX2 Inst_REgIDst_do_reg_11_ ( .D(n2644), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[11]) );
  SDFFRQX2 Inst_REgIDst_do_reg_12_ ( .D(n2646), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[12]) );
  SDFFRQX2 Inst_REgIDst_do_reg_13_ ( .D(n2648), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[13]) );
  SDFFRQX2 Inst_REgIDst_do_reg_14_ ( .D(n2650), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[14]) );
  SDFFRQX2 Inst_REgIDst_do_reg_15_ ( .D(n2652), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[15]) );
  SDFFRQX2 Inst_REgIDst_do_reg_16_ ( .D(n2654), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[16]) );
  SDFFRQX2 Inst_REgIDst_do_reg_17_ ( .D(n2656), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[17]) );
  SDFFRQX2 Inst_REgIDst_do_reg_18_ ( .D(n2658), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[18]) );
  SDFFRQX2 Inst_REgIDst_do_reg_19_ ( .D(n2660), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n170), .Q(IDstReg[19]) );
  SDFFRQX2 Inst_REgIDst_do_reg_20_ ( .D(n2662), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[20]) );
  SDFFRQX2 Inst_REgIDst_do_reg_21_ ( .D(n2664), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[21]) );
  SDFFRQX2 Inst_REgIDst_do_reg_22_ ( .D(n2666), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[22]) );
  SDFFRQX2 Inst_REgIDst_do_reg_23_ ( .D(n2668), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[23]) );
  SDFFRQX2 Inst_REgIDst_do_reg_24_ ( .D(n2670), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[24]) );
  SDFFRQX2 Inst_REgIDst_do_reg_25_ ( .D(n2672), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[25]) );
  SDFFRQX2 Inst_REgIDst_do_reg_26_ ( .D(n2674), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[26]) );
  SDFFRQX2 Inst_REgIDst_do_reg_27_ ( .D(n2676), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[27]) );
  SDFFRQX2 Inst_REgIDst_do_reg_28_ ( .D(n2678), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[28]) );
  SDFFRQX2 Inst_REgIDst_do_reg_29_ ( .D(n2680), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[29]) );
  SDFFRQX2 Inst_REgIDst_do_reg_30_ ( .D(n2682), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[30]) );
  SDFFRQX2 Inst_REgIDst_do_reg_31_ ( .D(n2684), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n171), .Q(IDstReg[31]) );
  SDFFRQX2 Inst_REgIDst_do_reg_32_ ( .D(n2686), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[32]) );
  SDFFRQX2 Inst_REgIDst_do_reg_33_ ( .D(n2688), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[33]) );
  SDFFRQX2 Inst_REgIDst_do_reg_34_ ( .D(n2690), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[34]) );
  SDFFRQX2 Inst_REgIDst_do_reg_35_ ( .D(n2692), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[35]) );
  SDFFRQX2 Inst_REgIDst_do_reg_36_ ( .D(n2694), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[36]) );
  SDFFRQX2 Inst_REgIDst_do_reg_37_ ( .D(n2696), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[37]) );
  SDFFRQX2 Inst_REgIDst_do_reg_38_ ( .D(n2698), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[38]) );
  SDFFRQX2 Inst_REgIDst_do_reg_39_ ( .D(n2700), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[39]) );
  SDFFRQX2 Inst_REgIDst_do_reg_40_ ( .D(n2702), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[40]) );
  SDFFRQX2 Inst_REgIDst_do_reg_41_ ( .D(n2704), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[41]) );
  SDFFRQX2 Inst_REgIDst_do_reg_42_ ( .D(n2706), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[42]) );
  SDFFRQX2 Inst_REgIDst_do_reg_43_ ( .D(n2708), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n172), .Q(IDstReg[43]) );
  SDFFRQX2 Inst_REgIDst_do_reg_44_ ( .D(n2710), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[44]) );
  SDFFRQX2 Inst_REgIDst_do_reg_45_ ( .D(n2712), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[45]) );
  SDFFRQX2 Inst_REgIDst_do_reg_46_ ( .D(n2714), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[46]) );
  SDFFRQX2 Inst_REgIDst_do_reg_47_ ( .D(n2716), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[47]) );
  SDFFRQX2 Inst_REgIDst_do_reg_48_ ( .D(n2718), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[48]) );
  SDFFRQX2 Inst_REgIDst_do_reg_49_ ( .D(n2720), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[49]) );
  SDFFRQX2 Inst_REgIDst_do_reg_50_ ( .D(n2722), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[50]) );
  SDFFRQX2 Inst_REgIDst_do_reg_51_ ( .D(n2724), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[51]) );
  SDFFRQX2 Inst_REgIDst_do_reg_52_ ( .D(n2726), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[52]) );
  SDFFRQX2 Inst_REgIDst_do_reg_53_ ( .D(n2728), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[53]) );
  SDFFRQX2 Inst_REgIDst_do_reg_54_ ( .D(n2730), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[54]) );
  SDFFRQX2 Inst_REgIDst_do_reg_55_ ( .D(n2732), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n173), .Q(IDstReg[55]) );
  SDFFRQX2 Inst_REgIDst_do_reg_56_ ( .D(n2734), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[56]) );
  SDFFRQX2 Inst_REgIDst_do_reg_57_ ( .D(n2736), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[57]) );
  SDFFRQX2 Inst_REgIDst_do_reg_58_ ( .D(n2738), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[58]) );
  SDFFRQX2 Inst_REgIDst_do_reg_59_ ( .D(n2740), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[59]) );
  SDFFRQX2 Inst_REgIDst_do_reg_60_ ( .D(n2742), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[60]) );
  SDFFRQX2 Inst_REgIDst_do_reg_61_ ( .D(n2744), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[61]) );
  SDFFRQX2 Inst_REgIDst_do_reg_62_ ( .D(n2746), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[62]) );
  SDFFRQX2 Inst_REgIDst_do_reg_63_ ( .D(n2748), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(n174), .Q(IDstReg[63]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_5_ ( .D(Inst_forkAE_REG_TK2_N7), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[101]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_17_ ( .D(Inst_forkAE_REG_TK2_N19), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[113]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_21_ ( .D(Inst_forkAE_REG_TK2_N23), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[117]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_25_ ( .D(Inst_forkAE_REG_TK2_N27), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[121]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_29_ ( .D(Inst_forkAE_REG_TK2_N31), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[125]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_48_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N50), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[48]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_52_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N54), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[52]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_60_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N62), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[60]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_16_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N18), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[16]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_20_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N22), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[20]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_28_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N30), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[28]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_56_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N58), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[56]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_24_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N26), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[24]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_2_ ( .D(Inst_forkAE_KEY_INVERSE[162]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[162]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_25_ ( .D(Inst_forkAE_KEY_INVERSE[185]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[185]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_29_ ( .D(Inst_forkAE_KEY_INVERSE[189]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[189]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_33_ ( .D(Inst_forkAE_KEY_INVERSE[145]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[145]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_34_ ( .D(Inst_forkAE_KEY_INVERSE[146]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[146]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_37_ ( .D(Inst_forkAE_KEY_INVERSE[141]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[141]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_38_ ( .D(Inst_forkAE_KEY_INVERSE[142]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[142]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_42_ ( .D(Inst_forkAE_KEY_INVERSE[134]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[134]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_3_ ( .D(Inst_forkAE_KEY_INVERSE[163]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[163]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_7_ ( .D(Inst_forkAE_KEY_INVERSE[167]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[167]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_9_ ( .D(Inst_forkAE_KEY_INVERSE[169]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[169]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_10_ ( .D(Inst_forkAE_KEY_INVERSE[170]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[170]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_13_ ( .D(Inst_forkAE_KEY_INVERSE[173]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[173]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_15_ ( .D(Inst_forkAE_KEY_INVERSE[175]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[175]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_19_ ( .D(Inst_forkAE_KEY_INVERSE[179]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[179]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_23_ ( .D(Inst_forkAE_KEY_INVERSE[183]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[183]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_27_ ( .D(Inst_forkAE_KEY_INVERSE[187]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[187]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_31_ ( .D(Inst_forkAE_KEY_INVERSE[191]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[191]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_32_ ( .D(Inst_forkAE_KEY_INVERSE[144]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[144]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_35_ ( .D(Inst_forkAE_KEY_INVERSE[147]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[147]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_39_ ( .D(Inst_forkAE_KEY_INVERSE[143]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[143]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_40_ ( .D(Inst_forkAE_KEY_INVERSE[132]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[132]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_43_ ( .D(Inst_forkAE_KEY_INVERSE[135]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[135]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_47_ ( .D(Inst_forkAE_KEY_INVERSE[151]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[151]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_0_ ( .D(Inst_forkAE_KEY_INVERSE[160]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[160]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_1_ ( .D(Inst_forkAE_KEY_INVERSE[161]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[161]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_4_ ( .D(Inst_forkAE_KEY_INVERSE[164]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[164]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_5_ ( .D(Inst_forkAE_KEY_INVERSE[165]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[165]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_6_ ( .D(Inst_forkAE_KEY_INVERSE[166]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[166]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_8_ ( .D(Inst_forkAE_KEY_INVERSE[168]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[168]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_11_ ( .D(Inst_forkAE_KEY_INVERSE[171]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[171]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_12_ ( .D(Inst_forkAE_KEY_INVERSE[172]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[172]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_14_ ( .D(Inst_forkAE_KEY_INVERSE[174]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[174]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_16_ ( .D(Inst_forkAE_KEY_INVERSE[176]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[176]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_17_ ( .D(Inst_forkAE_KEY_INVERSE[177]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[177]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_18_ ( .D(Inst_forkAE_KEY_INVERSE[178]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[178]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_20_ ( .D(Inst_forkAE_KEY_INVERSE[180]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[180]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_21_ ( .D(Inst_forkAE_KEY_INVERSE[181]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[181]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_22_ ( .D(Inst_forkAE_KEY_INVERSE[182]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[182]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_24_ ( .D(Inst_forkAE_KEY_INVERSE[184]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[184]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_26_ ( .D(Inst_forkAE_KEY_INVERSE[186]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[186]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_28_ ( .D(Inst_forkAE_KEY_INVERSE[188]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[188]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_30_ ( .D(Inst_forkAE_KEY_INVERSE[190]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[190]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_36_ ( .D(Inst_forkAE_KEY_INVERSE[140]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[140]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_53_ ( .D(Inst_forkAE_KEY_INVERSE[157]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[157]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_3_ ( .D(Inst_forkAE_L_N5), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[3]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_37_ ( .D(Inst_forkAE_L_N39), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[37]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_1_ ( .D(Inst_forkAE_L_N3), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[1]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_5_ ( .D(Inst_forkAE_L_N7), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[5]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_8_ ( .D(Inst_forkAE_L_N10), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(C1[8]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_32_ ( .D(Inst_forkAE_L_N34), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[32]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_14_ ( .D(Inst_forkAE_REG_TK2_0_N16), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[46]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_18_ ( .D(Inst_forkAE_REG_TK2_0_N20), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[50]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_26_ ( .D(Inst_forkAE_REG_TK2_0_N28), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[58]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_0_ ( .D(Inst_forkAE_REG_TK2_N2), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[96]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_28_ ( .D(Inst_forkAE_L_N30), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[28]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_10_ ( .D(Inst_forkAE_REG_TK2_0_N12), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[42]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_33_ ( .D(Inst_forkAE_REG_TK2_0_N35), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[18]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_34_ ( .D(Inst_forkAE_REG_TK2_0_N36), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[19]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_37_ ( .D(Inst_forkAE_REG_TK2_0_N39), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[14]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_38_ ( .D(Inst_forkAE_REG_TK2_0_N40), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[15]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_23_ ( .D(Inst_forkAE_L_N25), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[23]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_31_ ( .D(Inst_forkAE_L_N33), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[31]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_63_ ( .D(Inst_forkAE_L_N65), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[63]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_63_ ( .D(Inst_lfsr_n132), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[63]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_47_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N49), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[47]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_0_ ( .D(Inst_forkAE_L_N2), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[0]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_16_ ( .D(Inst_forkAE_L_N18), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[16]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_20_ ( .D(Inst_forkAE_L_N22), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[20]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_24_ ( .D(Inst_forkAE_L_N26), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[24]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_36_ ( .D(Inst_forkAE_L_N38), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[36]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_44_ ( .D(Inst_forkAE_L_N46), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[44]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_48_ ( .D(Inst_forkAE_L_N50), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[48]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_60_ ( .D(Inst_forkAE_L_N62), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[60]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_37_ ( .D(Inst_forkAE_REG_TK2_N39), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[76])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_57_ ( .D(Inst_forkAE_REG_TK2_N59), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[64])
         );
  SDFFSQXL Inst_forkAE_L_Q_reg_52_ ( .D(Inst_forkAE_L_N54), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[52]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_56_ ( .D(Inst_forkAE_L_N58), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[56]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_53_ ( .D(Inst_forkAE_REG_TK2_N55), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[92])
         );
  SDFFRQX2 Inst_RegIDt_do_reg_7_ ( .D(Inst_RegIDt_n17), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[7]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_8_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N10), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[8]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_19_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N21), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[19]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_23_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N25), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[23]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_27_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N29), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[27]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_31_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N33), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[31]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_32_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N34), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[32]) );
  SDFFRQX2 Inst_RegIDt_do_reg_0_ ( .D(Inst_RegIDt_n3), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[0]) );
  SDFFRQX2 Inst_RegIDt_do_reg_1_ ( .D(Inst_RegIDt_n5), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[1]) );
  SDFFRQX2 Inst_RegIDt_do_reg_2_ ( .D(Inst_RegIDt_n7), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[2]) );
  SDFFRQX2 Inst_RegIDt_do_reg_3_ ( .D(Inst_RegIDt_n9), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[3]) );
  SDFFRQX2 Inst_RegIDt_do_reg_4_ ( .D(Inst_RegIDt_n11), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[4]) );
  SDFFRQX2 Inst_RegIDt_do_reg_5_ ( .D(Inst_RegIDt_n13), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[5]) );
  SDFFRQX2 Inst_RegIDt_do_reg_6_ ( .D(Inst_RegIDt_n15), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[6]) );
  SDFFRQX2 Inst_RegIDt_do_reg_8_ ( .D(Inst_RegIDt_n19), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[8]) );
  SDFFRQX2 Inst_RegIDt_do_reg_9_ ( .D(Inst_RegIDt_n21), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[9]) );
  SDFFRQX2 Inst_RegIDt_do_reg_10_ ( .D(Inst_RegIDt_n23), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[10]) );
  SDFFRQX2 Inst_RegIDt_do_reg_11_ ( .D(Inst_RegIDt_n25), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n164), .Q(IDtReg[11]) );
  SDFFRQX2 Inst_RegIDt_do_reg_12_ ( .D(Inst_RegIDt_n27), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[12]) );
  SDFFRQX2 Inst_RegIDt_do_reg_13_ ( .D(Inst_RegIDt_n29), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[13]) );
  SDFFRQX2 Inst_RegIDt_do_reg_14_ ( .D(Inst_RegIDt_n31), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[14]) );
  SDFFRQX2 Inst_RegIDt_do_reg_15_ ( .D(Inst_RegIDt_n33), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[15]) );
  SDFFRQX2 Inst_RegIDt_do_reg_16_ ( .D(Inst_RegIDt_n35), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[16]) );
  SDFFRQX2 Inst_RegIDt_do_reg_17_ ( .D(Inst_RegIDt_n37), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[17]) );
  SDFFRQX2 Inst_RegIDt_do_reg_18_ ( .D(Inst_RegIDt_n39), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[18]) );
  SDFFRQX2 Inst_RegIDt_do_reg_19_ ( .D(Inst_RegIDt_n41), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[19]) );
  SDFFRQX2 Inst_RegIDt_do_reg_20_ ( .D(Inst_RegIDt_n43), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[20]) );
  SDFFRQX2 Inst_RegIDt_do_reg_21_ ( .D(Inst_RegIDt_n45), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[21]) );
  SDFFRQX2 Inst_RegIDt_do_reg_22_ ( .D(Inst_RegIDt_n47), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[22]) );
  SDFFRQX2 Inst_RegIDt_do_reg_23_ ( .D(Inst_RegIDt_n49), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n165), .Q(IDtReg[23]) );
  SDFFRQX2 Inst_RegIDt_do_reg_24_ ( .D(Inst_RegIDt_n51), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[24]) );
  SDFFRQX2 Inst_RegIDt_do_reg_25_ ( .D(Inst_RegIDt_n53), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[25]) );
  SDFFRQX2 Inst_RegIDt_do_reg_26_ ( .D(Inst_RegIDt_n55), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[26]) );
  SDFFRQX2 Inst_RegIDt_do_reg_27_ ( .D(Inst_RegIDt_n57), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[27]) );
  SDFFRQX2 Inst_RegIDt_do_reg_28_ ( .D(Inst_RegIDt_n59), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[28]) );
  SDFFRQX2 Inst_RegIDt_do_reg_29_ ( .D(Inst_RegIDt_n61), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[29]) );
  SDFFRQX2 Inst_RegIDt_do_reg_30_ ( .D(Inst_RegIDt_n63), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[30]) );
  SDFFRQX2 Inst_RegIDt_do_reg_31_ ( .D(Inst_RegIDt_n65), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[31]) );
  SDFFRQX2 Inst_RegIDt_do_reg_32_ ( .D(Inst_RegIDt_n67), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[32]) );
  SDFFRQX2 Inst_RegIDt_do_reg_33_ ( .D(Inst_RegIDt_n69), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[33]) );
  SDFFRQX2 Inst_RegIDt_do_reg_34_ ( .D(Inst_RegIDt_n71), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[34]) );
  SDFFRQX2 Inst_RegIDt_do_reg_35_ ( .D(Inst_RegIDt_n73), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n166), .Q(IDtReg[35]) );
  SDFFRQX2 Inst_RegIDt_do_reg_36_ ( .D(Inst_RegIDt_n75), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[36]) );
  SDFFRQX2 Inst_RegIDt_do_reg_37_ ( .D(Inst_RegIDt_n77), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[37]) );
  SDFFRQX2 Inst_RegIDt_do_reg_38_ ( .D(Inst_RegIDt_n79), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[38]) );
  SDFFRQX2 Inst_RegIDt_do_reg_39_ ( .D(Inst_RegIDt_n81), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[39]) );
  SDFFRQX2 Inst_RegIDt_do_reg_40_ ( .D(Inst_RegIDt_n83), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[40]) );
  SDFFRQX2 Inst_RegIDt_do_reg_41_ ( .D(Inst_RegIDt_n85), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[41]) );
  SDFFRQX2 Inst_RegIDt_do_reg_42_ ( .D(Inst_RegIDt_n87), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[42]) );
  SDFFRQX2 Inst_RegIDt_do_reg_43_ ( .D(Inst_RegIDt_n89), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[43]) );
  SDFFRQX2 Inst_RegIDt_do_reg_44_ ( .D(Inst_RegIDt_n91), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[44]) );
  SDFFRQX2 Inst_RegIDt_do_reg_45_ ( .D(Inst_RegIDt_n93), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[45]) );
  SDFFRQX2 Inst_RegIDt_do_reg_46_ ( .D(Inst_RegIDt_n95), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[46]) );
  SDFFRQX2 Inst_RegIDt_do_reg_47_ ( .D(Inst_RegIDt_n97), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n167), .Q(IDtReg[47]) );
  SDFFRQX2 Inst_RegIDt_do_reg_48_ ( .D(Inst_RegIDt_n99), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[48]) );
  SDFFRQX2 Inst_RegIDt_do_reg_49_ ( .D(Inst_RegIDt_n101), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[49]) );
  SDFFRQX2 Inst_RegIDt_do_reg_50_ ( .D(Inst_RegIDt_n103), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[50]) );
  SDFFRQX2 Inst_RegIDt_do_reg_51_ ( .D(Inst_RegIDt_n105), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[51]) );
  SDFFRQX2 Inst_RegIDt_do_reg_52_ ( .D(Inst_RegIDt_n107), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[52]) );
  SDFFRQX2 Inst_RegIDt_do_reg_53_ ( .D(Inst_RegIDt_n109), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[53]) );
  SDFFRQX2 Inst_RegIDt_do_reg_54_ ( .D(Inst_RegIDt_n111), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[54]) );
  SDFFRQX2 Inst_RegIDt_do_reg_55_ ( .D(Inst_RegIDt_n113), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[55]) );
  SDFFRQX2 Inst_RegIDt_do_reg_56_ ( .D(Inst_RegIDt_n115), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[56]) );
  SDFFRQX2 Inst_RegIDt_do_reg_57_ ( .D(Inst_RegIDt_n117), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[57]) );
  SDFFRQX2 Inst_RegIDt_do_reg_58_ ( .D(Inst_RegIDt_n119), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[58]) );
  SDFFRQX2 Inst_RegIDt_do_reg_59_ ( .D(Inst_RegIDt_n121), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n168), .Q(IDtReg[59]) );
  SDFFRQX2 Inst_RegIDt_do_reg_60_ ( .D(Inst_RegIDt_n123), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n169), .Q(IDtReg[60]) );
  SDFFRQX2 Inst_RegIDt_do_reg_61_ ( .D(Inst_RegIDt_n125), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n169), .Q(IDtReg[61]) );
  SDFFRQX2 Inst_RegIDt_do_reg_62_ ( .D(Inst_RegIDt_n127), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n169), .Q(IDtReg[62]) );
  SDFFRQX2 Inst_RegIDt_do_reg_63_ ( .D(Inst_RegIDt_n130), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .RN(n169), .Q(IDtReg[63]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_51_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N53), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[51]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_55_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N57), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[55]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_59_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N61), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[59]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_63_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N65), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[63]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_4_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N6), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[4]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_36_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N38), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[36]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_40_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N42), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[40]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_44_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N46), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[44]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_0_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N2), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[0]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_12_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N14), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[12]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_63_ ( .D(Inst_forkAE_KEY_INVERSE[155]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[155]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_44_ ( .D(Inst_forkAE_KEY_INVERSE[148]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[148]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_45_ ( .D(Inst_forkAE_KEY_INVERSE[149]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[149]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_46_ ( .D(Inst_forkAE_KEY_INVERSE[150]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[150]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_62_ ( .D(Inst_forkAE_KEY_INVERSE[154]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[154]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_2_ ( .D(Inst_forkAE_REG_TK2_0_N4), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[34])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_6_ ( .D(Inst_forkAE_REG_TK2_0_N8), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[38])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_22_ ( .D(Inst_forkAE_REG_TK2_0_N24), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[54]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_30_ ( .D(Inst_forkAE_REG_TK2_0_N32), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[62]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_50_ ( .D(Inst_forkAE_KEY_INVERSE[138]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[138]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_51_ ( .D(Inst_forkAE_KEY_INVERSE[139]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[139]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_55_ ( .D(Inst_forkAE_KEY_INVERSE[159]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[159]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_58_ ( .D(Inst_forkAE_KEY_INVERSE[130]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[130]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_59_ ( .D(Inst_forkAE_KEY_INVERSE[131]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[131]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_41_ ( .D(Inst_forkAE_KEY_INVERSE[133]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[133]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_54_ ( .D(Inst_forkAE_KEY_INVERSE[158]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[158]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_48_ ( .D(Inst_forkAE_KEY_INVERSE[136]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[136]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_49_ ( .D(Inst_forkAE_KEY_INVERSE[137]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[137]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_52_ ( .D(Inst_forkAE_KEY_INVERSE[156]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[156]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_56_ ( .D(Inst_forkAE_KEY_INVERSE[128]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[128]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_57_ ( .D(Inst_forkAE_KEY_INVERSE[129]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[129]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_60_ ( .D(Inst_forkAE_KEY_INVERSE[152]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[152]) );
  SDFFSQXL Inst_forkAE_REG_TK1_Q_reg_61_ ( .D(Inst_forkAE_KEY_INVERSE[153]), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[153]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_6_ ( .D(Inst_forkAE_L_N8), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[6]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_34_ ( .D(Inst_forkAE_L_N36), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[34]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_28_ ( .D(Inst_forkAE_REG_TK2_N30), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[124]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_8_ ( .D(Inst_forkAE_REG_TK2_N10), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[104]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_9_ ( .D(Inst_forkAE_L_N11), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(C1[9]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_2_ ( .D(Inst_forkAE_L_N4), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[2]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_21_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N23), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[21]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_29_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N31), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[29]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_10_ ( .D(Inst_forkAE_REG_TK2_N12), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[106]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_43_ ( .D(Inst_forkAE_L_N45), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[43]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_47_ ( .D(Inst_forkAE_L_N49), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[47]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_17_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N19), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[17]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_53_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N55), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[53]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_57_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N59), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[57]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_33_ ( .D(Inst_forkAE_REG_TK2_N35), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[80])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_45_ ( .D(Inst_forkAE_REG_TK2_N47), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[84])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_49_ ( .D(Inst_forkAE_REG_TK2_N51), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[72])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_61_ ( .D(Inst_forkAE_REG_TK2_N63), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[88])
         );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_25_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N27), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[25]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_49_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N51), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[49]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_61_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N63), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[61]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_41_ ( .D(Inst_forkAE_REG_TK2_N43), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[68])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_1_ ( .D(Inst_forkAE_REG_TK2_0_N3), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[33])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_41_ ( .D(Inst_forkAE_REG_TK2_0_N43), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[6]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_42_ ( .D(Inst_forkAE_REG_TK2_0_N44), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[7]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_12_ ( .D(Inst_forkAE_REG_TK2_N14), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[108]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_29_ ( .D(Inst_forkAE_L_N31), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[29]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_53_ ( .D(Inst_forkAE_L_N55), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[53]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_19_ ( .D(Inst_forkAE_L_N21), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[19]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_39_ ( .D(Inst_forkAE_L_N41), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[39]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_11_ ( .D(Inst_forkAE_L_N13), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[11]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_42_ ( .D(Inst_forkAE_REG_TK2_N44), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[69])
         );
  SDFFSQXL Inst_forkAE_L_Q_reg_49_ ( .D(Inst_forkAE_L_N51), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[49]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_61_ ( .D(Inst_forkAE_L_N63), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[61]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_55_ ( .D(Inst_forkAE_L_N57), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[55]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_59_ ( .D(Inst_forkAE_L_N61), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[59]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_5_ ( .D(Inst_forkAE_REG_TK2_0_N7), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[37])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_9_ ( .D(Inst_forkAE_REG_TK2_0_N11), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[41]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_13_ ( .D(Inst_forkAE_REG_TK2_0_N15), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[45]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_17_ ( .D(Inst_forkAE_REG_TK2_0_N19), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[49]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_21_ ( .D(Inst_forkAE_REG_TK2_0_N23), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[53]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_25_ ( .D(Inst_forkAE_REG_TK2_0_N27), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[57]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_29_ ( .D(Inst_forkAE_REG_TK2_0_N31), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[61]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_45_ ( .D(Inst_forkAE_REG_TK2_0_N47), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[22]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_46_ ( .D(Inst_forkAE_REG_TK2_0_N48), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[23]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_49_ ( .D(Inst_forkAE_REG_TK2_0_N51), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[10]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_50_ ( .D(Inst_forkAE_REG_TK2_0_N52), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[11]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_54_ ( .D(Inst_forkAE_REG_TK2_0_N56), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[31]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_57_ ( .D(Inst_forkAE_REG_TK2_0_N59), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[2]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_58_ ( .D(Inst_forkAE_REG_TK2_0_N60), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[3]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_61_ ( .D(Inst_forkAE_REG_TK2_0_N63), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[26]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_62_ ( .D(Inst_forkAE_REG_TK2_0_N64), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[27]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_2_ ( .D(Inst_forkAE_REG_TK2_N4), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[98]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_3_ ( .D(Inst_forkAE_REG_TK2_N5), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[99]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_14_ ( .D(Inst_forkAE_REG_TK2_N16), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[110]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_27_ ( .D(Inst_forkAE_L_N29), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[27]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_35_ ( .D(Inst_forkAE_L_N37), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[35]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_51_ ( .D(Inst_forkAE_L_N53), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[51]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_7_ ( .D(Inst_forkAE_L_N9), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(C1[7]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_38_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N40), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[38]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_50_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N52), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[50]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_58_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N60), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[58]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_1_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N3), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[1]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_3_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N5), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[3]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_5_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N7), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[5]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_7_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N9), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[7]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_13_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N15), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[13]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_43_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N45), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[43]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_15_ ( .D(Inst_forkAE_L_N17), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[15]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_18_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N20), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[18]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_26_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N28), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[26]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_30_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N32), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[30]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_22_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N24), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[22]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_54_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N56), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[54]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_62_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N64), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[62]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_35_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N37), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[35]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_39_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N41), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[39]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_11_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N13), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[11]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_15_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N17), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[15]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_4_ ( .D(Inst_forkAE_REG_TK2_N6), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[100]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_16_ ( .D(Inst_forkAE_REG_TK2_N18), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[112]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_20_ ( .D(Inst_forkAE_REG_TK2_N22), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[116]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_24_ ( .D(Inst_forkAE_REG_TK2_N26), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[120]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_25_ ( .D(Inst_forkAE_L_N27), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[25]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_57_ ( .D(Inst_forkAE_L_N59), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[57]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_13_ ( .D(Inst_forkAE_L_N15), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[13]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_33_ ( .D(Inst_forkAE_L_N35), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[33]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_41_ ( .D(Inst_forkAE_L_N43), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[41]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_53_ ( .D(Inst_forkAE_REG_TK2_0_N55), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[30]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_45_ ( .D(Inst_forkAE_L_N47), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[45]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_17_ ( .D(Inst_forkAE_L_N19), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[17]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_21_ ( .D(Inst_forkAE_L_N23), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[21]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_46_ ( .D(Inst_forkAE_L_N48), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[46]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_44_ ( .D(Inst_forkAE_REG_TK2_N46), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_108_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_52_ ( .D(Inst_forkAE_REG_TK2_N54), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_116_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_56_ ( .D(Inst_forkAE_REG_TK2_N58), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_120_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_60_ ( .D(Inst_forkAE_REG_TK2_N62), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_124_) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_33_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N35), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[33]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_55_ ( .D(Inst_forkAE_REG_TK2_N57), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[94])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_59_ ( .D(Inst_forkAE_REG_TK2_N61), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[66])
         );
  SDFFSQXL Inst_forkAE_L_Q_reg_26_ ( .D(Inst_forkAE_L_N28), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[26]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_50_ ( .D(Inst_forkAE_L_N52), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[50]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_9_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N11), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[9]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_18_ ( .D(Inst_forkAE_L_N20), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[18]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_22_ ( .D(Inst_forkAE_L_N24), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[22]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_11_ ( .D(Inst_forkAE_REG_TK2_N13), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[107]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_15_ ( .D(Inst_forkAE_REG_TK2_N17), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[111]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_58_ ( .D(Inst_forkAE_L_N60), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[58]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_62_ ( .D(Inst_forkAE_L_N64), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[62]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_37_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N39), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[37]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_41_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N43), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[41]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_0_ ( .D(Inst_forkAE_REG_TK2_0_N2), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[32])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_47_ ( .D(Inst_forkAE_REG_TK2_0_N49), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_47_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_34_ ( .D(Inst_forkAE_REG_TK2_N36), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[81])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_38_ ( .D(Inst_forkAE_REG_TK2_N40), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[77])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_39_ ( .D(Inst_forkAE_REG_TK2_N41), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[78])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_46_ ( .D(Inst_forkAE_REG_TK2_N48), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[85])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_50_ ( .D(Inst_forkAE_REG_TK2_N52), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[73])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_54_ ( .D(Inst_forkAE_REG_TK2_N56), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[93])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_58_ ( .D(Inst_forkAE_REG_TK2_N60), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[65])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_62_ ( .D(Inst_forkAE_REG_TK2_N64), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[89])
         );
  SDFFSQXL Inst_forkAE_L_Q_reg_30_ ( .D(Inst_forkAE_L_N32), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[30]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_54_ ( .D(Inst_forkAE_L_N56), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[54]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_14_ ( .D(Inst_forkAE_L_N16), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[14]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_42_ ( .D(Inst_forkAE_L_N44), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[42]) );
  SDFFSQXL Inst_forkAE_FSM_X_state_reg_1_ ( .D(Inst_forkAE_FSM_X_N42), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_FSM_X_state_1_)
         );
  SDFFSQXL Inst_forkAE_L_Q_reg_10_ ( .D(Inst_forkAE_L_N12), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[10]) );
  SDFFSQXL Inst_forkAE_L_Q_reg_38_ ( .D(Inst_forkAE_L_N40), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(C1[38]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_32_ ( .D(Inst_forkAE_REG_TK2_N34), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_96_)
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_36_ ( .D(Inst_forkAE_REG_TK2_N38), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_100_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_40_ ( .D(Inst_forkAE_REG_TK2_N42), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_104_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_48_ ( .D(Inst_forkAE_REG_TK2_N50), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CURRENT_KEY_112_) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_42_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N44), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[42]) );
  SDFFSQXL Inst_forkAE_ConstGen_STATE_reg_6_ ( .D(Inst_forkAE_ConstGen_N30), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CONST_DEC_6_) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_1_ ( .D(Inst_forkAE_REG_TK2_N3), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[97]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_13_ ( .D(Inst_forkAE_REG_TK2_N15), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[109]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_34_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N36), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[34]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_6_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N8), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[6]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_9_ ( .D(Inst_forkAE_REG_TK2_N11), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[105]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_10_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N12), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[10]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_46_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N48), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[46]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_0_ ( .D(Inst_lfsr_n195), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[0]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_45_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N47), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[45]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_2_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N4), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[2]) );
  SDFFSQXL Inst_forkAE_REG_INTERNAL_STATE_Q_reg_14_ ( .D(
        Inst_forkAE_REG_INTERNAL_STATE_N16), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .SN(1'b1), .Q(C0[14]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_51_ ( .D(Inst_forkAE_REG_TK2_N53), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[74])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_63_ ( .D(Inst_forkAE_REG_TK2_N65), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[90])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_11_ ( .D(Inst_forkAE_REG_TK2_0_N13), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[43]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_7_ ( .D(Inst_forkAE_REG_TK2_N9), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[103]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_23_ ( .D(Inst_forkAE_REG_TK2_N25), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[119]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_47_ ( .D(Inst_forkAE_REG_TK2_N49), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[86])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_3_ ( .D(Inst_forkAE_REG_TK2_0_N5), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[35])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_7_ ( .D(Inst_forkAE_REG_TK2_0_N9), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[39])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_23_ ( .D(Inst_forkAE_REG_TK2_0_N25), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[55]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_31_ ( .D(Inst_forkAE_REG_TK2_0_N33), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[63]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_6_ ( .D(Inst_forkAE_REG_TK2_N8), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[102]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_22_ ( .D(Inst_forkAE_REG_TK2_N24), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[118]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_31_ ( .D(Inst_forkAE_REG_TK2_N33), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[127]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_36_ ( .D(Inst_forkAE_REG_TK2_0_N38), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[13]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_44_ ( .D(Inst_forkAE_REG_TK2_0_N46), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[21]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_48_ ( .D(Inst_forkAE_REG_TK2_0_N50), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[9]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_52_ ( .D(Inst_forkAE_REG_TK2_0_N54), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[29]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_56_ ( .D(Inst_forkAE_REG_TK2_0_N58), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[1]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_60_ ( .D(Inst_forkAE_REG_TK2_0_N62), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[25]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_27_ ( .D(Inst_forkAE_REG_TK2_N29), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[123]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_32_ ( .D(Inst_forkAE_REG_TK2_0_N34), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[17]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_40_ ( .D(Inst_forkAE_REG_TK2_0_N42), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[5]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_19_ ( .D(Inst_forkAE_REG_TK2_N21), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[115]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_35_ ( .D(Inst_forkAE_REG_TK2_N37), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[82])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_43_ ( .D(Inst_forkAE_REG_TK2_N45), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[70])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_35_ ( .D(Inst_forkAE_REG_TK2_0_N37), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_35_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_39_ ( .D(Inst_forkAE_REG_TK2_0_N41), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_39_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_43_ ( .D(Inst_forkAE_REG_TK2_0_N45), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_43_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_55_ ( .D(Inst_forkAE_REG_TK2_0_N57), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_55_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_59_ ( .D(Inst_forkAE_REG_TK2_0_N61), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_59_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_63_ ( .D(Inst_forkAE_REG_TK2_0_N65), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_63_) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_15_ ( .D(Inst_forkAE_REG_TK2_0_N17), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[47]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_19_ ( .D(Inst_forkAE_REG_TK2_0_N21), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[51]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_27_ ( .D(Inst_forkAE_REG_TK2_0_N29), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[59]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_18_ ( .D(Inst_forkAE_REG_TK2_N20), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[114]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_26_ ( .D(Inst_forkAE_REG_TK2_N28), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[122]) );
  SDFFSQXL Inst_forkAE_REG_TK2_Q_reg_30_ ( .D(Inst_forkAE_REG_TK2_N32), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[126]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_8_ ( .D(Inst_forkAE_REG_TK2_0_N10), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[40]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_4_ ( .D(Inst_forkAE_REG_TK2_0_N6), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_KEY_INVERSE[36])
         );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_12_ ( .D(Inst_forkAE_REG_TK2_0_N14), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[44]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_16_ ( .D(Inst_forkAE_REG_TK2_0_N18), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[48]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_20_ ( .D(Inst_forkAE_REG_TK2_0_N22), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[52]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_24_ ( .D(Inst_forkAE_REG_TK2_0_N26), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[56]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_28_ ( .D(Inst_forkAE_REG_TK2_0_N30), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_KEY_INVERSE[60]) );
  SDFFSQXL Inst_forkAE_REG_TK2_0_Q_reg_51_ ( .D(Inst_forkAE_REG_TK2_0_N53), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(
        Inst_forkAE_CURRENT_KEY_51_) );
  SDFFSQXL Inst_forkAE_FSM_X_state_reg_2_ ( .D(Inst_forkAE_FSM_X_N43), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_FSM_X_state_2_)
         );
  SDFFSQXL Inst_forkAE_ConstGen_STATE_reg_4_ ( .D(Inst_forkAE_ConstGen_N28), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CONST_ENC_5_) );
  SDFFSQXL Inst_lfsr_counter_up_reg_62_ ( .D(Inst_lfsr_n133), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[62]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_61_ ( .D(Inst_lfsr_n134), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[61]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_59_ ( .D(Inst_lfsr_n136), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[59]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_58_ ( .D(Inst_lfsr_n137), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[58]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_57_ ( .D(Inst_lfsr_n138), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[57]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_55_ ( .D(Inst_lfsr_n140), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[55]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_54_ ( .D(Inst_lfsr_n141), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[54]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_53_ ( .D(Inst_lfsr_n142), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[53]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_51_ ( .D(Inst_lfsr_n144), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[51]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_50_ ( .D(Inst_lfsr_n145), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[50]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_49_ ( .D(Inst_lfsr_n146), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[49]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_47_ ( .D(Inst_lfsr_n148), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[47]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_46_ ( .D(Inst_lfsr_n149), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[46]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_45_ ( .D(Inst_lfsr_n150), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[45]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_43_ ( .D(Inst_lfsr_n152), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[43]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_42_ ( .D(Inst_lfsr_n153), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[42]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_41_ ( .D(Inst_lfsr_n154), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[41]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_39_ ( .D(Inst_lfsr_n156), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[39]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_38_ ( .D(Inst_lfsr_n157), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[38]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_37_ ( .D(Inst_lfsr_n158), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[37]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_35_ ( .D(Inst_lfsr_n160), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[35]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_34_ ( .D(Inst_lfsr_n161), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[34]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_33_ ( .D(Inst_lfsr_n162), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[33]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_31_ ( .D(Inst_lfsr_n164), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[31]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_30_ ( .D(Inst_lfsr_n165), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[30]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_29_ ( .D(Inst_lfsr_n166), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[29]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_28_ ( .D(Inst_lfsr_n167), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[28]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_27_ ( .D(Inst_lfsr_n168), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[27]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_26_ ( .D(Inst_lfsr_n169), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[26]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_25_ ( .D(Inst_lfsr_n170), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[25]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_24_ ( .D(Inst_lfsr_n171), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[24]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_23_ ( .D(Inst_lfsr_n172), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[23]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_22_ ( .D(Inst_lfsr_n173), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[22]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_21_ ( .D(Inst_lfsr_n174), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[21]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_20_ ( .D(Inst_lfsr_n175), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[20]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_19_ ( .D(Inst_lfsr_n176), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[19]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_18_ ( .D(Inst_lfsr_n177), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[18]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_17_ ( .D(Inst_lfsr_n178), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[17]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_16_ ( .D(Inst_lfsr_n179), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[16]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_15_ ( .D(Inst_lfsr_n180), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[15]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_14_ ( .D(Inst_lfsr_n181), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[14]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_13_ ( .D(Inst_lfsr_n182), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[13]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_12_ ( .D(Inst_lfsr_n183), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[12]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_11_ ( .D(Inst_lfsr_n184), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[11]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_10_ ( .D(Inst_lfsr_n185), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[10]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_9_ ( .D(Inst_lfsr_n186), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[9]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_8_ ( .D(Inst_lfsr_n187), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[8]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_7_ ( .D(Inst_lfsr_n188), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[7]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_6_ ( .D(Inst_lfsr_n189), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[6]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_5_ ( .D(Inst_lfsr_n190), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[5]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_4_ ( .D(Inst_lfsr_n191), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[4]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_3_ ( .D(Inst_lfsr_n192), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[3]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_2_ ( .D(Inst_lfsr_n193), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[2]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_1_ ( .D(Inst_lfsr_n194), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[1]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_60_ ( .D(Inst_lfsr_n135), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[60]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_56_ ( .D(Inst_lfsr_n139), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[56]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_52_ ( .D(Inst_lfsr_n143), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[52]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_48_ ( .D(Inst_lfsr_n147), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[48]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_44_ ( .D(Inst_lfsr_n151), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[44]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_40_ ( .D(Inst_lfsr_n155), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[40]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_36_ ( .D(Inst_lfsr_n159), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[36]) );
  SDFFSQXL Inst_lfsr_counter_up_reg_32_ ( .D(Inst_lfsr_n163), .SI(1'b0), .SE(
        1'b0), .CK(clk), .SN(1'b1), .Q(randd[32]) );
  SDFFSQXL Inst_forkAE_FSM_X_state_reg_0_ ( .D(Inst_forkAE_FSM_X_N41), .SI(
        1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_FSM_X_state_0_)
         );
  SDFFSQXL Inst_forkAE_ConstGen_STATE_reg_1_ ( .D(Inst_forkAE_ConstGen_N25), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CONST_ENC_2_) );
  SDFFSQXL Inst_forkAE_ConstGen_STATE_reg_0_ ( .D(Inst_forkAE_ConstGen_N24), 
        .SI(1'b0), .SE(1'b0), .CK(clk), .SN(1'b1), .Q(Inst_forkAE_CONST_ENC_1_) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_62 ( .A(randd[62]), .B(
        Inst_lfsr_add_3205_carry[62]), .CO(Inst_lfsr_add_3205_carry[63]), .S(
        Inst_lfsr_N66) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_61 ( .A(randd[61]), .B(
        Inst_lfsr_add_3205_carry[61]), .CO(Inst_lfsr_add_3205_carry[62]), .S(
        Inst_lfsr_N65) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_60 ( .A(randd[60]), .B(
        Inst_lfsr_add_3205_carry[60]), .CO(Inst_lfsr_add_3205_carry[61]), .S(
        Inst_lfsr_N64) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_59 ( .A(randd[59]), .B(
        Inst_lfsr_add_3205_carry[59]), .CO(Inst_lfsr_add_3205_carry[60]), .S(
        Inst_lfsr_N63) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_58 ( .A(randd[58]), .B(
        Inst_lfsr_add_3205_carry[58]), .CO(Inst_lfsr_add_3205_carry[59]), .S(
        Inst_lfsr_N62) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_57 ( .A(randd[57]), .B(
        Inst_lfsr_add_3205_carry[57]), .CO(Inst_lfsr_add_3205_carry[58]), .S(
        Inst_lfsr_N61) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_56 ( .A(randd[56]), .B(
        Inst_lfsr_add_3205_carry[56]), .CO(Inst_lfsr_add_3205_carry[57]), .S(
        Inst_lfsr_N60) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_55 ( .A(randd[55]), .B(
        Inst_lfsr_add_3205_carry[55]), .CO(Inst_lfsr_add_3205_carry[56]), .S(
        Inst_lfsr_N59) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_54 ( .A(randd[54]), .B(
        Inst_lfsr_add_3205_carry[54]), .CO(Inst_lfsr_add_3205_carry[55]), .S(
        Inst_lfsr_N58) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_53 ( .A(randd[53]), .B(
        Inst_lfsr_add_3205_carry[53]), .CO(Inst_lfsr_add_3205_carry[54]), .S(
        Inst_lfsr_N57) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_52 ( .A(randd[52]), .B(
        Inst_lfsr_add_3205_carry[52]), .CO(Inst_lfsr_add_3205_carry[53]), .S(
        Inst_lfsr_N56) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_51 ( .A(randd[51]), .B(
        Inst_lfsr_add_3205_carry[51]), .CO(Inst_lfsr_add_3205_carry[52]), .S(
        Inst_lfsr_N55) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_50 ( .A(randd[50]), .B(
        Inst_lfsr_add_3205_carry[50]), .CO(Inst_lfsr_add_3205_carry[51]), .S(
        Inst_lfsr_N54) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_49 ( .A(randd[49]), .B(
        Inst_lfsr_add_3205_carry[49]), .CO(Inst_lfsr_add_3205_carry[50]), .S(
        Inst_lfsr_N53) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_48 ( .A(randd[48]), .B(
        Inst_lfsr_add_3205_carry[48]), .CO(Inst_lfsr_add_3205_carry[49]), .S(
        Inst_lfsr_N52) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_47 ( .A(randd[47]), .B(
        Inst_lfsr_add_3205_carry[47]), .CO(Inst_lfsr_add_3205_carry[48]), .S(
        Inst_lfsr_N51) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_46 ( .A(randd[46]), .B(
        Inst_lfsr_add_3205_carry[46]), .CO(Inst_lfsr_add_3205_carry[47]), .S(
        Inst_lfsr_N50) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_45 ( .A(randd[45]), .B(
        Inst_lfsr_add_3205_carry[45]), .CO(Inst_lfsr_add_3205_carry[46]), .S(
        Inst_lfsr_N49) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_44 ( .A(randd[44]), .B(
        Inst_lfsr_add_3205_carry[44]), .CO(Inst_lfsr_add_3205_carry[45]), .S(
        Inst_lfsr_N48) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_43 ( .A(randd[43]), .B(
        Inst_lfsr_add_3205_carry[43]), .CO(Inst_lfsr_add_3205_carry[44]), .S(
        Inst_lfsr_N47) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_42 ( .A(randd[42]), .B(
        Inst_lfsr_add_3205_carry[42]), .CO(Inst_lfsr_add_3205_carry[43]), .S(
        Inst_lfsr_N46) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_41 ( .A(randd[41]), .B(
        Inst_lfsr_add_3205_carry[41]), .CO(Inst_lfsr_add_3205_carry[42]), .S(
        Inst_lfsr_N45) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_40 ( .A(randd[40]), .B(
        Inst_lfsr_add_3205_carry[40]), .CO(Inst_lfsr_add_3205_carry[41]), .S(
        Inst_lfsr_N44) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_39 ( .A(randd[39]), .B(
        Inst_lfsr_add_3205_carry[39]), .CO(Inst_lfsr_add_3205_carry[40]), .S(
        Inst_lfsr_N43) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_38 ( .A(randd[38]), .B(
        Inst_lfsr_add_3205_carry[38]), .CO(Inst_lfsr_add_3205_carry[39]), .S(
        Inst_lfsr_N42) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_37 ( .A(randd[37]), .B(
        Inst_lfsr_add_3205_carry[37]), .CO(Inst_lfsr_add_3205_carry[38]), .S(
        Inst_lfsr_N41) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_36 ( .A(randd[36]), .B(
        Inst_lfsr_add_3205_carry[36]), .CO(Inst_lfsr_add_3205_carry[37]), .S(
        Inst_lfsr_N40) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_35 ( .A(randd[35]), .B(
        Inst_lfsr_add_3205_carry[35]), .CO(Inst_lfsr_add_3205_carry[36]), .S(
        Inst_lfsr_N39) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_34 ( .A(randd[34]), .B(
        Inst_lfsr_add_3205_carry[34]), .CO(Inst_lfsr_add_3205_carry[35]), .S(
        Inst_lfsr_N38) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_33 ( .A(randd[33]), .B(
        Inst_lfsr_add_3205_carry[33]), .CO(Inst_lfsr_add_3205_carry[34]), .S(
        Inst_lfsr_N37) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_32 ( .A(randd[32]), .B(
        Inst_lfsr_add_3205_carry[32]), .CO(Inst_lfsr_add_3205_carry[33]), .S(
        Inst_lfsr_N36) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_31 ( .A(randd[31]), .B(
        Inst_lfsr_add_3205_carry[31]), .CO(Inst_lfsr_add_3205_carry[32]), .S(
        Inst_lfsr_N35) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_30 ( .A(randd[30]), .B(
        Inst_lfsr_add_3205_carry[30]), .CO(Inst_lfsr_add_3205_carry[31]), .S(
        Inst_lfsr_N34) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_29 ( .A(randd[29]), .B(
        Inst_lfsr_add_3205_carry[29]), .CO(Inst_lfsr_add_3205_carry[30]), .S(
        Inst_lfsr_N33) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_28 ( .A(randd[28]), .B(
        Inst_lfsr_add_3205_carry[28]), .CO(Inst_lfsr_add_3205_carry[29]), .S(
        Inst_lfsr_N32) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_27 ( .A(randd[27]), .B(
        Inst_lfsr_add_3205_carry[27]), .CO(Inst_lfsr_add_3205_carry[28]), .S(
        Inst_lfsr_N31) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_26 ( .A(randd[26]), .B(
        Inst_lfsr_add_3205_carry[26]), .CO(Inst_lfsr_add_3205_carry[27]), .S(
        Inst_lfsr_N30) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_25 ( .A(randd[25]), .B(
        Inst_lfsr_add_3205_carry[25]), .CO(Inst_lfsr_add_3205_carry[26]), .S(
        Inst_lfsr_N29) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_24 ( .A(randd[24]), .B(
        Inst_lfsr_add_3205_carry[24]), .CO(Inst_lfsr_add_3205_carry[25]), .S(
        Inst_lfsr_N28) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_23 ( .A(randd[23]), .B(
        Inst_lfsr_add_3205_carry[23]), .CO(Inst_lfsr_add_3205_carry[24]), .S(
        Inst_lfsr_N27) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_22 ( .A(randd[22]), .B(
        Inst_lfsr_add_3205_carry[22]), .CO(Inst_lfsr_add_3205_carry[23]), .S(
        Inst_lfsr_N26) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_21 ( .A(randd[21]), .B(
        Inst_lfsr_add_3205_carry[21]), .CO(Inst_lfsr_add_3205_carry[22]), .S(
        Inst_lfsr_N25) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_20 ( .A(randd[20]), .B(
        Inst_lfsr_add_3205_carry[20]), .CO(Inst_lfsr_add_3205_carry[21]), .S(
        Inst_lfsr_N24) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_19 ( .A(randd[19]), .B(
        Inst_lfsr_add_3205_carry[19]), .CO(Inst_lfsr_add_3205_carry[20]), .S(
        Inst_lfsr_N23) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_18 ( .A(randd[18]), .B(
        Inst_lfsr_add_3205_carry[18]), .CO(Inst_lfsr_add_3205_carry[19]), .S(
        Inst_lfsr_N22) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_17 ( .A(randd[17]), .B(
        Inst_lfsr_add_3205_carry[17]), .CO(Inst_lfsr_add_3205_carry[18]), .S(
        Inst_lfsr_N21) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_16 ( .A(randd[16]), .B(
        Inst_lfsr_add_3205_carry[16]), .CO(Inst_lfsr_add_3205_carry[17]), .S(
        Inst_lfsr_N20) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_15 ( .A(randd[15]), .B(
        Inst_lfsr_add_3205_carry[15]), .CO(Inst_lfsr_add_3205_carry[16]), .S(
        Inst_lfsr_N19) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_14 ( .A(randd[14]), .B(
        Inst_lfsr_add_3205_carry[14]), .CO(Inst_lfsr_add_3205_carry[15]), .S(
        Inst_lfsr_N18) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_13 ( .A(randd[13]), .B(
        Inst_lfsr_add_3205_carry[13]), .CO(Inst_lfsr_add_3205_carry[14]), .S(
        Inst_lfsr_N17) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_12 ( .A(randd[12]), .B(
        Inst_lfsr_add_3205_carry[12]), .CO(Inst_lfsr_add_3205_carry[13]), .S(
        Inst_lfsr_N16) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_11 ( .A(randd[11]), .B(
        Inst_lfsr_add_3205_carry[11]), .CO(Inst_lfsr_add_3205_carry[12]), .S(
        Inst_lfsr_N15) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_10 ( .A(randd[10]), .B(
        Inst_lfsr_add_3205_carry[10]), .CO(Inst_lfsr_add_3205_carry[11]), .S(
        Inst_lfsr_N14) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_9 ( .A(randd[9]), .B(
        Inst_lfsr_add_3205_carry[9]), .CO(Inst_lfsr_add_3205_carry[10]), .S(
        Inst_lfsr_N13) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_8 ( .A(randd[8]), .B(
        Inst_lfsr_add_3205_carry[8]), .CO(Inst_lfsr_add_3205_carry[9]), .S(
        Inst_lfsr_N12) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_7 ( .A(randd[7]), .B(
        Inst_lfsr_add_3205_carry[7]), .CO(Inst_lfsr_add_3205_carry[8]), .S(
        Inst_lfsr_N11) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_6 ( .A(randd[6]), .B(
        Inst_lfsr_add_3205_carry[6]), .CO(Inst_lfsr_add_3205_carry[7]), .S(
        Inst_lfsr_N10) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_5 ( .A(randd[5]), .B(
        Inst_lfsr_add_3205_carry[5]), .CO(Inst_lfsr_add_3205_carry[6]), .S(
        Inst_lfsr_N9) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_4 ( .A(randd[4]), .B(
        Inst_lfsr_add_3205_carry[4]), .CO(Inst_lfsr_add_3205_carry[5]), .S(
        Inst_lfsr_N8) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_3 ( .A(randd[3]), .B(
        Inst_lfsr_add_3205_carry[3]), .CO(Inst_lfsr_add_3205_carry[4]), .S(
        Inst_lfsr_N7) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_2 ( .A(randd[2]), .B(
        Inst_lfsr_add_3205_carry[2]), .CO(Inst_lfsr_add_3205_carry[3]), .S(
        Inst_lfsr_N6) );
  ADDHX1 Inst_lfsr_add_3205_U1_1_1 ( .A(randd[1]), .B(randd[0]), .CO(
        Inst_lfsr_add_3205_carry[2]), .S(Inst_lfsr_N5) );
  OR2X2 U259 ( .A(n135), .B(n184), .Y(n1245) );
  OR2X2 U260 ( .A(n1242), .B(n964), .Y(n961) );
  NOR2X2 U261 ( .A(n187), .B(rst), .Y(n186) );
  NOR2X4 U262 ( .A(rst), .B(en_c), .Y(n187) );
  NOR3X6 U263 ( .A(n963), .B(n1243), .C(n184), .Y(n964) );
  INVX2 U264 ( .A(n1244), .Y(n963) );
  INVXL U265 ( .A(n1251), .Y(n134) );
  INVX2 U266 ( .A(n134), .Y(n135) );
  AND3X4 U267 ( .A(n944), .B(n945), .C(n145), .Y(n210) );
  INVX2 U268 ( .A(n1249), .Y(n1257) );
  NOR3X8 U269 ( .A(n136), .B(n944), .C(n945), .Y(n196) );
  CLKINVX3 U270 ( .A(n233), .Y(n193) );
  NAND3X2 U271 ( .A(n145), .B(n944), .C(n947), .Y(n233) );
  BUFX2 U272 ( .A(n162), .Y(n153) );
  BUFX2 U273 ( .A(n160), .Y(n158) );
  BUFX2 U274 ( .A(n161), .Y(n154) );
  BUFX2 U275 ( .A(n161), .Y(n155) );
  BUFX2 U276 ( .A(n161), .Y(n156) );
  BUFX2 U277 ( .A(n160), .Y(n157) );
  BUFX2 U278 ( .A(n162), .Y(n151) );
  BUFX2 U279 ( .A(n162), .Y(n152) );
  BUFX2 U280 ( .A(n160), .Y(n159) );
  BUFX2 U281 ( .A(n194), .Y(n160) );
  BUFX2 U282 ( .A(n194), .Y(n161) );
  BUFX2 U283 ( .A(n194), .Y(n162) );
  BUFX2 U284 ( .A(n175), .Y(n173) );
  BUFX2 U285 ( .A(n175), .Y(n172) );
  BUFX2 U286 ( .A(n176), .Y(n171) );
  BUFX2 U287 ( .A(n176), .Y(n170) );
  BUFX2 U288 ( .A(n176), .Y(n169) );
  BUFX2 U289 ( .A(n177), .Y(n168) );
  BUFX2 U290 ( .A(n177), .Y(n167) );
  BUFX2 U291 ( .A(n177), .Y(n166) );
  BUFX2 U292 ( .A(n178), .Y(n165) );
  BUFX2 U293 ( .A(n178), .Y(n164) );
  BUFX2 U294 ( .A(n175), .Y(n174) );
  BUFX2 U295 ( .A(n148), .Y(n138) );
  BUFX2 U296 ( .A(n148), .Y(n139) );
  BUFX2 U297 ( .A(n146), .Y(n144) );
  BUFX2 U298 ( .A(n147), .Y(n143) );
  BUFX2 U299 ( .A(n146), .Y(n145) );
  BUFX2 U300 ( .A(n147), .Y(n141) );
  BUFX2 U301 ( .A(n148), .Y(n140) );
  BUFX2 U302 ( .A(n147), .Y(n142) );
  BUFX2 U303 ( .A(n163), .Y(n150) );
  BUFX2 U304 ( .A(n194), .Y(n163) );
  INVX2 U305 ( .A(n146), .Y(n136) );
  BUFX2 U306 ( .A(n2105), .Y(n175) );
  BUFX2 U307 ( .A(n2105), .Y(n176) );
  BUFX2 U308 ( .A(n2105), .Y(n177) );
  BUFX2 U309 ( .A(n2105), .Y(n178) );
  BUFX2 U310 ( .A(n190), .Y(n146) );
  BUFX2 U311 ( .A(n190), .Y(n148) );
  BUFX2 U312 ( .A(n190), .Y(n147) );
  BUFX2 U313 ( .A(n149), .Y(n137) );
  BUFX2 U314 ( .A(n190), .Y(n149) );
  CLKINVX1 U315 ( .A(rst), .Y(n2105) );
  MXI2X1 U316 ( .A(n182), .B(n183), .S0(n184), .Y(n2106) );
  MXI2X1 U317 ( .A(n183), .B(n179), .S0(n184), .Y(n2107) );
  MXI2X1 U318 ( .A(n180), .B(n185), .S0(n184), .Y(n2108) );
  MX2X1 U319 ( .A(n186), .B(n187), .S0(randd[0]), .Y(Inst_lfsr_n195) );
  AO22X1 U320 ( .A0(n187), .A1(randd[1]), .B0(Inst_lfsr_N5), .B1(n186), .Y(
        Inst_lfsr_n194) );
  AO22X1 U321 ( .A0(n187), .A1(randd[2]), .B0(Inst_lfsr_N6), .B1(n186), .Y(
        Inst_lfsr_n193) );
  AO22X1 U322 ( .A0(n187), .A1(randd[3]), .B0(Inst_lfsr_N7), .B1(n186), .Y(
        Inst_lfsr_n192) );
  AO22X1 U323 ( .A0(n187), .A1(randd[4]), .B0(Inst_lfsr_N8), .B1(n186), .Y(
        Inst_lfsr_n191) );
  AO22X1 U324 ( .A0(n187), .A1(randd[5]), .B0(Inst_lfsr_N9), .B1(n186), .Y(
        Inst_lfsr_n190) );
  AO22X1 U325 ( .A0(n187), .A1(randd[6]), .B0(Inst_lfsr_N10), .B1(n186), .Y(
        Inst_lfsr_n189) );
  AO22X1 U326 ( .A0(n187), .A1(randd[7]), .B0(Inst_lfsr_N11), .B1(n186), .Y(
        Inst_lfsr_n188) );
  AO22X1 U327 ( .A0(n187), .A1(randd[8]), .B0(Inst_lfsr_N12), .B1(n186), .Y(
        Inst_lfsr_n187) );
  AO22X1 U328 ( .A0(n187), .A1(randd[9]), .B0(Inst_lfsr_N13), .B1(n186), .Y(
        Inst_lfsr_n186) );
  AO22X1 U329 ( .A0(n187), .A1(randd[10]), .B0(Inst_lfsr_N14), .B1(n186), .Y(
        Inst_lfsr_n185) );
  AO22X1 U330 ( .A0(n187), .A1(randd[11]), .B0(Inst_lfsr_N15), .B1(n186), .Y(
        Inst_lfsr_n184) );
  AO22X1 U331 ( .A0(n187), .A1(randd[12]), .B0(Inst_lfsr_N16), .B1(n186), .Y(
        Inst_lfsr_n183) );
  AO22X1 U332 ( .A0(n187), .A1(randd[13]), .B0(Inst_lfsr_N17), .B1(n186), .Y(
        Inst_lfsr_n182) );
  AO22X1 U333 ( .A0(n187), .A1(randd[14]), .B0(Inst_lfsr_N18), .B1(n186), .Y(
        Inst_lfsr_n181) );
  AO22X1 U334 ( .A0(n187), .A1(randd[15]), .B0(Inst_lfsr_N19), .B1(n186), .Y(
        Inst_lfsr_n180) );
  AO22X1 U335 ( .A0(n187), .A1(randd[16]), .B0(Inst_lfsr_N20), .B1(n186), .Y(
        Inst_lfsr_n179) );
  AO22X1 U336 ( .A0(n187), .A1(randd[17]), .B0(Inst_lfsr_N21), .B1(n186), .Y(
        Inst_lfsr_n178) );
  AO22X1 U337 ( .A0(n187), .A1(randd[18]), .B0(Inst_lfsr_N22), .B1(n186), .Y(
        Inst_lfsr_n177) );
  AO22X1 U338 ( .A0(n187), .A1(randd[19]), .B0(Inst_lfsr_N23), .B1(n186), .Y(
        Inst_lfsr_n176) );
  AO22X1 U339 ( .A0(n187), .A1(randd[20]), .B0(Inst_lfsr_N24), .B1(n186), .Y(
        Inst_lfsr_n175) );
  AO22X1 U340 ( .A0(n187), .A1(randd[21]), .B0(Inst_lfsr_N25), .B1(n186), .Y(
        Inst_lfsr_n174) );
  AO22X1 U341 ( .A0(n187), .A1(randd[22]), .B0(Inst_lfsr_N26), .B1(n186), .Y(
        Inst_lfsr_n173) );
  AO22X1 U342 ( .A0(n187), .A1(randd[23]), .B0(Inst_lfsr_N27), .B1(n186), .Y(
        Inst_lfsr_n172) );
  AO22X1 U343 ( .A0(n187), .A1(randd[24]), .B0(Inst_lfsr_N28), .B1(n186), .Y(
        Inst_lfsr_n171) );
  AO22X1 U344 ( .A0(n187), .A1(randd[25]), .B0(Inst_lfsr_N29), .B1(n186), .Y(
        Inst_lfsr_n170) );
  AO22X1 U345 ( .A0(n187), .A1(randd[26]), .B0(Inst_lfsr_N30), .B1(n186), .Y(
        Inst_lfsr_n169) );
  AO22X1 U346 ( .A0(n187), .A1(randd[27]), .B0(Inst_lfsr_N31), .B1(n186), .Y(
        Inst_lfsr_n168) );
  AO22X1 U347 ( .A0(n187), .A1(randd[28]), .B0(Inst_lfsr_N32), .B1(n186), .Y(
        Inst_lfsr_n167) );
  AO22X1 U348 ( .A0(n187), .A1(randd[29]), .B0(Inst_lfsr_N33), .B1(n186), .Y(
        Inst_lfsr_n166) );
  AO22X1 U349 ( .A0(n187), .A1(randd[30]), .B0(Inst_lfsr_N34), .B1(n186), .Y(
        Inst_lfsr_n165) );
  AO22X1 U350 ( .A0(n187), .A1(randd[31]), .B0(Inst_lfsr_N35), .B1(n186), .Y(
        Inst_lfsr_n164) );
  AO22X1 U351 ( .A0(n187), .A1(randd[32]), .B0(Inst_lfsr_N36), .B1(n186), .Y(
        Inst_lfsr_n163) );
  AO22X1 U352 ( .A0(n187), .A1(randd[33]), .B0(Inst_lfsr_N37), .B1(n186), .Y(
        Inst_lfsr_n162) );
  AO22X1 U353 ( .A0(n187), .A1(randd[34]), .B0(Inst_lfsr_N38), .B1(n186), .Y(
        Inst_lfsr_n161) );
  AO22X1 U354 ( .A0(n187), .A1(randd[35]), .B0(Inst_lfsr_N39), .B1(n186), .Y(
        Inst_lfsr_n160) );
  AO22X1 U355 ( .A0(n187), .A1(randd[36]), .B0(Inst_lfsr_N40), .B1(n186), .Y(
        Inst_lfsr_n159) );
  AO22X1 U356 ( .A0(n187), .A1(randd[37]), .B0(Inst_lfsr_N41), .B1(n186), .Y(
        Inst_lfsr_n158) );
  AO22X1 U357 ( .A0(n187), .A1(randd[38]), .B0(Inst_lfsr_N42), .B1(n186), .Y(
        Inst_lfsr_n157) );
  AO22X1 U358 ( .A0(n187), .A1(randd[39]), .B0(Inst_lfsr_N43), .B1(n186), .Y(
        Inst_lfsr_n156) );
  AO22X1 U359 ( .A0(n187), .A1(randd[40]), .B0(Inst_lfsr_N44), .B1(n186), .Y(
        Inst_lfsr_n155) );
  AO22X1 U360 ( .A0(n187), .A1(randd[41]), .B0(Inst_lfsr_N45), .B1(n186), .Y(
        Inst_lfsr_n154) );
  AO22X1 U361 ( .A0(n187), .A1(randd[42]), .B0(Inst_lfsr_N46), .B1(n186), .Y(
        Inst_lfsr_n153) );
  AO22X1 U362 ( .A0(n187), .A1(randd[43]), .B0(Inst_lfsr_N47), .B1(n186), .Y(
        Inst_lfsr_n152) );
  AO22X1 U363 ( .A0(n187), .A1(randd[44]), .B0(Inst_lfsr_N48), .B1(n186), .Y(
        Inst_lfsr_n151) );
  AO22X1 U364 ( .A0(n187), .A1(randd[45]), .B0(Inst_lfsr_N49), .B1(n186), .Y(
        Inst_lfsr_n150) );
  AO22X1 U365 ( .A0(n187), .A1(randd[46]), .B0(Inst_lfsr_N50), .B1(n186), .Y(
        Inst_lfsr_n149) );
  AO22X1 U366 ( .A0(n187), .A1(randd[47]), .B0(Inst_lfsr_N51), .B1(n186), .Y(
        Inst_lfsr_n148) );
  AO22X1 U367 ( .A0(n187), .A1(randd[48]), .B0(Inst_lfsr_N52), .B1(n186), .Y(
        Inst_lfsr_n147) );
  AO22X1 U368 ( .A0(n187), .A1(randd[49]), .B0(Inst_lfsr_N53), .B1(n186), .Y(
        Inst_lfsr_n146) );
  AO22X1 U369 ( .A0(n187), .A1(randd[50]), .B0(Inst_lfsr_N54), .B1(n186), .Y(
        Inst_lfsr_n145) );
  AO22X1 U370 ( .A0(n187), .A1(randd[51]), .B0(Inst_lfsr_N55), .B1(n186), .Y(
        Inst_lfsr_n144) );
  AO22X1 U371 ( .A0(n187), .A1(randd[52]), .B0(Inst_lfsr_N56), .B1(n186), .Y(
        Inst_lfsr_n143) );
  AO22X1 U372 ( .A0(n187), .A1(randd[53]), .B0(Inst_lfsr_N57), .B1(n186), .Y(
        Inst_lfsr_n142) );
  AO22X1 U373 ( .A0(n187), .A1(randd[54]), .B0(Inst_lfsr_N58), .B1(n186), .Y(
        Inst_lfsr_n141) );
  AO22X1 U374 ( .A0(n187), .A1(randd[55]), .B0(Inst_lfsr_N59), .B1(n186), .Y(
        Inst_lfsr_n140) );
  AO22X1 U375 ( .A0(n187), .A1(randd[56]), .B0(Inst_lfsr_N60), .B1(n186), .Y(
        Inst_lfsr_n139) );
  AO22X1 U376 ( .A0(n187), .A1(randd[57]), .B0(Inst_lfsr_N61), .B1(n186), .Y(
        Inst_lfsr_n138) );
  AO22X1 U377 ( .A0(n187), .A1(randd[58]), .B0(Inst_lfsr_N62), .B1(n186), .Y(
        Inst_lfsr_n137) );
  AO22X1 U378 ( .A0(n187), .A1(randd[59]), .B0(Inst_lfsr_N63), .B1(n186), .Y(
        Inst_lfsr_n136) );
  AO22X1 U379 ( .A0(n187), .A1(randd[60]), .B0(Inst_lfsr_N64), .B1(n186), .Y(
        Inst_lfsr_n135) );
  AO22X1 U380 ( .A0(n187), .A1(randd[61]), .B0(Inst_lfsr_N65), .B1(n186), .Y(
        Inst_lfsr_n134) );
  AO22X1 U381 ( .A0(n187), .A1(randd[62]), .B0(Inst_lfsr_N66), .B1(n186), .Y(
        Inst_lfsr_n133) );
  MXI2X1 U382 ( .A(n188), .B(n189), .S0(randd[63]), .Y(Inst_lfsr_n132) );
  AOI2B1X1 U383 ( .A1N(Inst_lfsr_add_3205_carry[63]), .A0(n186), .B0(n187), 
        .Y(n189) );
  CLKNAND2X2 U384 ( .A(Inst_lfsr_add_3205_carry[63]), .B(n186), .Y(n188) );
  OAI2B11X1 U385 ( .A1N(Inst_forkAE_KEY_INVERSE[39]), .A0(n139), .B0(n191), 
        .C0(n192), .Y(Inst_forkAE_REG_TK2_0_N9) );
  AOI222XL U386 ( .A0(Inst_forkAE_KEY_INVERSE[7]), .A1(n193), .B0(n151), .B1(
        n195), .C0(n196), .C1(n197), .Y(n192) );
  MXI2X1 U387 ( .A(n198), .B(n199), .S0(Inst_forkAE_KEY_INVERSE[59]), .Y(n191)
         );
  OAI2B11X1 U388 ( .A1N(Inst_forkAE_KEY_INVERSE[38]), .A0(n137), .B0(n200), 
        .C0(n201), .Y(Inst_forkAE_REG_TK2_0_N8) );
  AOI222XL U389 ( .A0(Inst_forkAE_KEY_INVERSE[6]), .A1(n193), .B0(n150), .B1(
        n202), .C0(n196), .C1(n203), .Y(n201) );
  MXI2X1 U390 ( .A(n198), .B(n199), .S0(Inst_forkAE_KEY_INVERSE[56]), .Y(n200)
         );
  OAI211XL U391 ( .A0(n143), .A1(n204), .B0(n205), .C0(n206), .Y(
        Inst_forkAE_REG_TK2_0_N7) );
  AOI222XL U392 ( .A0(Inst_forkAE_KEY_INVERSE[5]), .A1(n193), .B0(n150), .B1(
        n207), .C0(n196), .C1(n208), .Y(n206) );
  MXI2X1 U393 ( .A(n198), .B(n199), .S0(n209), .Y(n205) );
  NOR2BX1 U394 ( .AN(n210), .B(n211), .Y(n199) );
  AND2X1 U395 ( .A(n210), .B(n211), .Y(n198) );
  OAI2B11X1 U396 ( .A1N(Inst_forkAE_CURRENT_KEY_63_), .A0(n137), .B0(n212), 
        .C0(n213), .Y(Inst_forkAE_REG_TK2_0_N65) );
  AOI222XL U397 ( .A0(Inst_forkAE_KEY_INVERSE[63]), .A1(n193), .B0(n196), .B1(
        n214), .C0(n154), .C1(n215), .Y(n213) );
  XOR2X1 U398 ( .A(n216), .B(n217), .Y(n214) );
  MXI2X1 U399 ( .A(n218), .B(n219), .S0(Inst_forkAE_CURRENT_KEY_43_), .Y(n212)
         );
  OAI211XL U400 ( .A0(n142), .A1(n220), .B0(n221), .C0(n222), .Y(
        Inst_forkAE_REG_TK2_0_N64) );
  AOI222XL U401 ( .A0(Inst_forkAE_KEY_INVERSE[62]), .A1(n193), .B0(n150), .B1(
        n223), .C0(n196), .C1(n216), .Y(n222) );
  MXI2X1 U402 ( .A(n218), .B(n219), .S0(Inst_forkAE_KEY_INVERSE[5]), .Y(n221)
         );
  OAI211XL U403 ( .A0(n143), .A1(n224), .B0(n225), .C0(n226), .Y(
        Inst_forkAE_REG_TK2_0_N63) );
  AOI222XL U404 ( .A0(Inst_forkAE_KEY_INVERSE[61]), .A1(n193), .B0(n150), .B1(
        n227), .C0(n196), .C1(n228), .Y(n226) );
  MXI2X1 U405 ( .A(n218), .B(n219), .S0(n229), .Y(n225) );
  NOR2BX1 U406 ( .AN(n210), .B(n230), .Y(n219) );
  AND2X1 U407 ( .A(n210), .B(n230), .Y(n218) );
  XOR2X1 U408 ( .A(n231), .B(n232), .Y(n230) );
  OAI221X1 U409 ( .A0(n233), .A1(n234), .B0(n139), .B1(n235), .C0(n236), .Y(
        Inst_forkAE_REG_TK2_0_N62) );
  AOI222XL U410 ( .A0(n196), .A1(n237), .B0(n210), .B1(n238), .C0(n154), .C1(
        n239), .Y(n236) );
  CLKINVX1 U411 ( .A(n240), .Y(n239) );
  XOR2X1 U412 ( .A(Inst_forkAE_KEY_INVERSE[6]), .B(n229), .Y(n238) );
  XOR2X1 U413 ( .A(Inst_forkAE_CURRENT_KEY_43_), .B(Inst_forkAE_KEY_INVERSE[5]), .Y(n229) );
  CLKINVX1 U414 ( .A(Inst_forkAE_KEY_INVERSE[25]), .Y(n235) );
  OAI2B11X1 U415 ( .A1N(Inst_forkAE_CURRENT_KEY_59_), .A0(n138), .B0(n241), 
        .C0(n242), .Y(Inst_forkAE_REG_TK2_0_N61) );
  AOI222XL U416 ( .A0(Inst_forkAE_KEY_INVERSE[59]), .A1(n193), .B0(n196), .B1(
        n243), .C0(n155), .C1(n244), .Y(n242) );
  XOR2X1 U417 ( .A(n245), .B(n246), .Y(n243) );
  MXI2X1 U418 ( .A(n247), .B(n248), .S0(Inst_forkAE_CURRENT_KEY_39_), .Y(n241)
         );
  OAI211XL U419 ( .A0(n143), .A1(n249), .B0(n250), .C0(n251), .Y(
        Inst_forkAE_REG_TK2_0_N60) );
  AOI222XL U420 ( .A0(Inst_forkAE_KEY_INVERSE[58]), .A1(n193), .B0(n150), .B1(
        n252), .C0(n196), .C1(n245), .Y(n251) );
  MXI2X1 U421 ( .A(n247), .B(n248), .S0(Inst_forkAE_KEY_INVERSE[13]), .Y(n250)
         );
  OAI221X1 U422 ( .A0(n253), .A1(n254), .B0(n140), .B1(n255), .C0(n256), .Y(
        Inst_forkAE_REG_TK2_0_N6) );
  AOI222XL U423 ( .A0(n153), .A1(n257), .B0(n193), .B1(n258), .C0(n210), .C1(
        n259), .Y(n256) );
  XOR2X1 U424 ( .A(Inst_forkAE_KEY_INVERSE[57]), .B(n209), .Y(n259) );
  XOR2X1 U425 ( .A(Inst_forkAE_KEY_INVERSE[59]), .B(
        Inst_forkAE_KEY_INVERSE[56]), .Y(n209) );
  XOR2X1 U426 ( .A(Inst_forkAE_KEY_INVERSE[7]), .B(Inst_forkAE_CURRENT_KEY_43_), .Y(n258) );
  OAI211XL U427 ( .A0(n142), .A1(n260), .B0(n261), .C0(n262), .Y(
        Inst_forkAE_REG_TK2_0_N59) );
  AOI222XL U428 ( .A0(Inst_forkAE_KEY_INVERSE[57]), .A1(n193), .B0(n150), .B1(
        n263), .C0(n196), .C1(n264), .Y(n262) );
  MXI2X1 U429 ( .A(n247), .B(n248), .S0(n265), .Y(n261) );
  NOR2BX1 U430 ( .AN(n210), .B(n266), .Y(n248) );
  AND2X1 U431 ( .A(n210), .B(n266), .Y(n247) );
  XOR2X1 U432 ( .A(n267), .B(n268), .Y(n266) );
  OAI221X1 U433 ( .A0(n233), .A1(n269), .B0(n140), .B1(n270), .C0(n271), .Y(
        Inst_forkAE_REG_TK2_0_N58) );
  AOI222XL U434 ( .A0(n196), .A1(n272), .B0(n210), .B1(n273), .C0(n154), .C1(
        n274), .Y(n271) );
  CLKINVX1 U435 ( .A(n275), .Y(n274) );
  XOR2X1 U436 ( .A(Inst_forkAE_KEY_INVERSE[14]), .B(n265), .Y(n273) );
  XOR2X1 U437 ( .A(Inst_forkAE_CURRENT_KEY_39_), .B(
        Inst_forkAE_KEY_INVERSE[13]), .Y(n265) );
  CLKINVX1 U438 ( .A(Inst_forkAE_KEY_INVERSE[1]), .Y(n270) );
  OAI2B11X1 U439 ( .A1N(Inst_forkAE_CURRENT_KEY_55_), .A0(n137), .B0(n276), 
        .C0(n277), .Y(Inst_forkAE_REG_TK2_0_N57) );
  AOI222XL U440 ( .A0(Inst_forkAE_KEY_INVERSE[55]), .A1(n193), .B0(n196), .B1(
        n278), .C0(n154), .C1(n279), .Y(n277) );
  XOR2X1 U441 ( .A(n280), .B(n281), .Y(n278) );
  MXI2X1 U442 ( .A(n282), .B(n283), .S0(Inst_forkAE_CURRENT_KEY_51_), .Y(n276)
         );
  OAI211XL U443 ( .A0(n142), .A1(n284), .B0(n285), .C0(n286), .Y(
        Inst_forkAE_REG_TK2_0_N56) );
  AOI222XL U444 ( .A0(Inst_forkAE_KEY_INVERSE[54]), .A1(n193), .B0(n150), .B1(
        n287), .C0(n196), .C1(n280), .Y(n286) );
  MXI2X1 U445 ( .A(n282), .B(n283), .S0(Inst_forkAE_KEY_INVERSE[9]), .Y(n285)
         );
  OAI2B11X1 U446 ( .A1N(Inst_forkAE_KEY_INVERSE[30]), .A0(n138), .B0(n288), 
        .C0(n289), .Y(Inst_forkAE_REG_TK2_0_N55) );
  AOI222XL U447 ( .A0(Inst_forkAE_KEY_INVERSE[53]), .A1(n193), .B0(n150), .B1(
        n290), .C0(n196), .C1(n291), .Y(n289) );
  MXI2X1 U448 ( .A(n282), .B(n283), .S0(n292), .Y(n288) );
  NOR2BX1 U449 ( .AN(n210), .B(n293), .Y(n283) );
  AND2X1 U450 ( .A(n210), .B(n293), .Y(n282) );
  XOR2X1 U451 ( .A(n294), .B(n295), .Y(n293) );
  OAI221X1 U452 ( .A0(n233), .A1(n296), .B0(n141), .B1(n297), .C0(n298), .Y(
        Inst_forkAE_REG_TK2_0_N54) );
  AOI222XL U453 ( .A0(n196), .A1(n299), .B0(n210), .B1(n300), .C0(n154), .C1(
        n301), .Y(n298) );
  CLKINVX1 U454 ( .A(n302), .Y(n301) );
  XOR2X1 U455 ( .A(Inst_forkAE_KEY_INVERSE[10]), .B(n292), .Y(n300) );
  XOR2X1 U456 ( .A(Inst_forkAE_CURRENT_KEY_51_), .B(Inst_forkAE_KEY_INVERSE[9]), .Y(n292) );
  CLKINVX1 U457 ( .A(Inst_forkAE_KEY_INVERSE[29]), .Y(n297) );
  OAI211XL U458 ( .A0(n142), .A1(n303), .B0(n304), .C0(n305), .Y(
        Inst_forkAE_REG_TK2_0_N53) );
  AOI222XL U459 ( .A0(Inst_forkAE_KEY_INVERSE[51]), .A1(n193), .B0(n196), .B1(
        n306), .C0(n155), .C1(n307), .Y(n305) );
  XOR2X1 U460 ( .A(n308), .B(n309), .Y(n306) );
  MXI2X1 U461 ( .A(n310), .B(n311), .S0(Inst_forkAE_CURRENT_KEY_55_), .Y(n304)
         );
  CLKINVX1 U462 ( .A(Inst_forkAE_CURRENT_KEY_51_), .Y(n303) );
  OAI211XL U463 ( .A0(n143), .A1(n295), .B0(n312), .C0(n313), .Y(
        Inst_forkAE_REG_TK2_0_N52) );
  AOI222XL U464 ( .A0(Inst_forkAE_KEY_INVERSE[50]), .A1(n193), .B0(n151), .B1(
        n314), .C0(n196), .C1(n308), .Y(n313) );
  MXI2X1 U465 ( .A(n310), .B(n311), .S0(Inst_forkAE_KEY_INVERSE[29]), .Y(n312)
         );
  CLKINVX1 U466 ( .A(Inst_forkAE_KEY_INVERSE[11]), .Y(n295) );
  OAI211XL U467 ( .A0(n143), .A1(n294), .B0(n315), .C0(n316), .Y(
        Inst_forkAE_REG_TK2_0_N51) );
  AOI222XL U468 ( .A0(Inst_forkAE_KEY_INVERSE[49]), .A1(n193), .B0(n150), .B1(
        n317), .C0(n196), .C1(n318), .Y(n316) );
  MXI2X1 U469 ( .A(n310), .B(n311), .S0(n319), .Y(n315) );
  NOR2BX1 U470 ( .AN(n210), .B(n320), .Y(n311) );
  AND2X1 U471 ( .A(n210), .B(n320), .Y(n310) );
  XNOR2X1 U472 ( .A(n284), .B(Inst_forkAE_KEY_INVERSE[30]), .Y(n320) );
  CLKINVX1 U473 ( .A(Inst_forkAE_KEY_INVERSE[31]), .Y(n284) );
  CLKINVX1 U474 ( .A(Inst_forkAE_KEY_INVERSE[10]), .Y(n294) );
  OAI221X1 U475 ( .A0(n233), .A1(n321), .B0(n141), .B1(n322), .C0(n323), .Y(
        Inst_forkAE_REG_TK2_0_N50) );
  AOI222XL U476 ( .A0(n196), .A1(n324), .B0(n210), .B1(n325), .C0(n154), .C1(
        n326), .Y(n323) );
  CLKINVX1 U477 ( .A(n327), .Y(n326) );
  XOR2X1 U478 ( .A(Inst_forkAE_KEY_INVERSE[30]), .B(n319), .Y(n325) );
  XOR2X1 U479 ( .A(Inst_forkAE_CURRENT_KEY_55_), .B(
        Inst_forkAE_KEY_INVERSE[29]), .Y(n319) );
  CLKINVX1 U480 ( .A(Inst_forkAE_KEY_INVERSE[9]), .Y(n322) );
  OAI2B11X1 U481 ( .A1N(Inst_forkAE_KEY_INVERSE[35]), .A0(n137), .B0(n328), 
        .C0(n329), .Y(Inst_forkAE_REG_TK2_0_N5) );
  AOI222XL U482 ( .A0(Inst_forkAE_KEY_INVERSE[3]), .A1(n193), .B0(n151), .B1(
        n245), .C0(n196), .C1(n330), .Y(n329) );
  XNOR2X1 U483 ( .A(n331), .B(randd[3]), .Y(n245) );
  CLKNAND2X2 U484 ( .A(IDtReg[3]), .B(MuxSel2), .Y(n331) );
  MXI2X1 U485 ( .A(n332), .B(n333), .S0(Inst_forkAE_KEY_INVERSE[47]), .Y(n328)
         );
  OAI211XL U486 ( .A0(n143), .A1(n334), .B0(n335), .C0(n336), .Y(
        Inst_forkAE_REG_TK2_0_N49) );
  AOI222XL U487 ( .A0(Inst_forkAE_KEY_INVERSE[47]), .A1(n193), .B0(n196), .B1(
        n337), .C0(n154), .C1(n338), .Y(n336) );
  XOR2X1 U488 ( .A(n339), .B(n340), .Y(n337) );
  MXI2X1 U489 ( .A(n341), .B(n342), .S0(Inst_forkAE_CURRENT_KEY_35_), .Y(n335)
         );
  OAI211XL U490 ( .A0(n142), .A1(n343), .B0(n344), .C0(n345), .Y(
        Inst_forkAE_REG_TK2_0_N48) );
  AOI222XL U491 ( .A0(Inst_forkAE_KEY_INVERSE[46]), .A1(n193), .B0(n151), .B1(
        n346), .C0(n196), .C1(n339), .Y(n345) );
  MXI2X1 U492 ( .A(n341), .B(n342), .S0(Inst_forkAE_KEY_INVERSE[17]), .Y(n344)
         );
  OAI211XL U493 ( .A0(n143), .A1(n347), .B0(n348), .C0(n349), .Y(
        Inst_forkAE_REG_TK2_0_N47) );
  AOI222XL U494 ( .A0(Inst_forkAE_KEY_INVERSE[45]), .A1(n193), .B0(n151), .B1(
        n350), .C0(n196), .C1(n351), .Y(n349) );
  MXI2X1 U495 ( .A(n341), .B(n342), .S0(n352), .Y(n348) );
  NOR2BX1 U496 ( .AN(n210), .B(n353), .Y(n342) );
  AND2X1 U497 ( .A(n210), .B(n353), .Y(n341) );
  XOR2X1 U498 ( .A(n354), .B(n355), .Y(n353) );
  OAI221X1 U499 ( .A0(n233), .A1(n356), .B0(n141), .B1(n357), .C0(n358), .Y(
        Inst_forkAE_REG_TK2_0_N46) );
  AOI222XL U500 ( .A0(n196), .A1(n359), .B0(n210), .B1(n360), .C0(n154), .C1(
        n361), .Y(n358) );
  CLKINVX1 U501 ( .A(n362), .Y(n361) );
  XOR2X1 U502 ( .A(Inst_forkAE_KEY_INVERSE[18]), .B(n352), .Y(n360) );
  XOR2X1 U503 ( .A(Inst_forkAE_CURRENT_KEY_35_), .B(
        Inst_forkAE_KEY_INVERSE[17]), .Y(n352) );
  CLKINVX1 U504 ( .A(Inst_forkAE_KEY_INVERSE[21]), .Y(n357) );
  OAI2B11X1 U505 ( .A1N(Inst_forkAE_CURRENT_KEY_43_), .A0(n138), .B0(n363), 
        .C0(n364), .Y(Inst_forkAE_REG_TK2_0_N45) );
  AOI222XL U506 ( .A0(Inst_forkAE_KEY_INVERSE[43]), .A1(n193), .B0(n196), .B1(
        n365), .C0(n155), .C1(n366), .Y(n364) );
  XOR2X1 U507 ( .A(n195), .B(n257), .Y(n365) );
  XNOR2X1 U508 ( .A(n367), .B(randd[4]), .Y(n257) );
  CLKNAND2X2 U509 ( .A(IDtReg[4]), .B(MuxSel2), .Y(n367) );
  MXI2X1 U510 ( .A(n368), .B(n369), .S0(Inst_forkAE_CURRENT_KEY_63_), .Y(n363)
         );
  OAI211XL U511 ( .A0(n232), .A1(n145), .B0(n370), .C0(n371), .Y(
        Inst_forkAE_REG_TK2_0_N44) );
  AOI222XL U512 ( .A0(Inst_forkAE_KEY_INVERSE[42]), .A1(n193), .B0(n151), .B1(
        n372), .C0(n196), .C1(n195), .Y(n371) );
  XNOR2X1 U513 ( .A(n373), .B(randd[7]), .Y(n195) );
  CLKNAND2X2 U514 ( .A(MuxSel2), .B(IDtReg[7]), .Y(n373) );
  MXI2X1 U515 ( .A(n368), .B(n369), .S0(Inst_forkAE_KEY_INVERSE[25]), .Y(n370)
         );
  CLKINVX1 U516 ( .A(Inst_forkAE_KEY_INVERSE[7]), .Y(n232) );
  OAI211XL U517 ( .A0(n143), .A1(n231), .B0(n374), .C0(n375), .Y(
        Inst_forkAE_REG_TK2_0_N43) );
  AOI222XL U518 ( .A0(Inst_forkAE_KEY_INVERSE[41]), .A1(n193), .B0(n151), .B1(
        n376), .C0(n196), .C1(n202), .Y(n375) );
  XNOR2X1 U519 ( .A(n377), .B(randd[6]), .Y(n202) );
  CLKNAND2X2 U520 ( .A(IDtReg[6]), .B(MuxSel2), .Y(n377) );
  MXI2X1 U521 ( .A(n368), .B(n369), .S0(n378), .Y(n374) );
  NOR2BX1 U522 ( .AN(n210), .B(n379), .Y(n369) );
  AND2X1 U523 ( .A(n210), .B(n379), .Y(n368) );
  XOR2X1 U524 ( .A(n224), .B(n220), .Y(n379) );
  CLKINVX1 U525 ( .A(Inst_forkAE_KEY_INVERSE[27]), .Y(n220) );
  CLKINVX1 U526 ( .A(Inst_forkAE_KEY_INVERSE[26]), .Y(n224) );
  CLKINVX1 U527 ( .A(Inst_forkAE_KEY_INVERSE[6]), .Y(n231) );
  OAI221X1 U528 ( .A0(n233), .A1(n380), .B0(n142), .B1(n381), .C0(n382), .Y(
        Inst_forkAE_REG_TK2_0_N42) );
  AOI222XL U529 ( .A0(n196), .A1(n207), .B0(n210), .B1(n383), .C0(n154), .C1(
        n384), .Y(n382) );
  CLKINVX1 U530 ( .A(n385), .Y(n384) );
  XOR2X1 U531 ( .A(Inst_forkAE_KEY_INVERSE[26]), .B(n378), .Y(n383) );
  XOR2X1 U532 ( .A(Inst_forkAE_CURRENT_KEY_63_), .B(
        Inst_forkAE_KEY_INVERSE[25]), .Y(n378) );
  XNOR2X1 U533 ( .A(n386), .B(randd[5]), .Y(n207) );
  CLKNAND2X2 U534 ( .A(IDtReg[5]), .B(MuxSel2), .Y(n386) );
  CLKINVX1 U535 ( .A(Inst_forkAE_KEY_INVERSE[5]), .Y(n381) );
  OAI2B11X1 U536 ( .A1N(Inst_forkAE_CURRENT_KEY_39_), .A0(n139), .B0(n387), 
        .C0(n388), .Y(Inst_forkAE_REG_TK2_0_N41) );
  AOI222XL U537 ( .A0(Inst_forkAE_KEY_INVERSE[39]), .A1(n193), .B0(n196), .B1(
        n389), .C0(n155), .C1(n197), .Y(n388) );
  XNOR2X1 U538 ( .A(n390), .B(randd[39]), .Y(n197) );
  CLKNAND2X2 U539 ( .A(IDtReg[39]), .B(MuxSel2), .Y(n390) );
  XOR2X1 U540 ( .A(n391), .B(n392), .Y(n389) );
  MXI2X1 U541 ( .A(n393), .B(n394), .S0(Inst_forkAE_CURRENT_KEY_59_), .Y(n387)
         );
  OAI211XL U542 ( .A0(n143), .A1(n268), .B0(n395), .C0(n396), .Y(
        Inst_forkAE_REG_TK2_0_N40) );
  AOI222XL U543 ( .A0(Inst_forkAE_KEY_INVERSE[38]), .A1(n193), .B0(n150), .B1(
        n203), .C0(n196), .C1(n391), .Y(n396) );
  XNOR2X1 U544 ( .A(n397), .B(randd[38]), .Y(n203) );
  CLKNAND2X2 U545 ( .A(IDtReg[38]), .B(MuxSel2), .Y(n397) );
  MXI2X1 U546 ( .A(n393), .B(n394), .S0(Inst_forkAE_KEY_INVERSE[1]), .Y(n395)
         );
  OAI2B11X1 U547 ( .A1N(Inst_forkAE_KEY_INVERSE[34]), .A0(n138), .B0(n398), 
        .C0(n399), .Y(Inst_forkAE_REG_TK2_0_N4) );
  AOI222XL U548 ( .A0(Inst_forkAE_KEY_INVERSE[2]), .A1(n193), .B0(n152), .B1(
        n264), .C0(n196), .C1(n400), .Y(n399) );
  XNOR2X1 U549 ( .A(n401), .B(randd[2]), .Y(n264) );
  CLKNAND2X2 U550 ( .A(IDtReg[2]), .B(MuxSel2), .Y(n401) );
  MXI2X1 U551 ( .A(n332), .B(n333), .S0(Inst_forkAE_KEY_INVERSE[44]), .Y(n398)
         );
  OAI211XL U552 ( .A0(n143), .A1(n267), .B0(n402), .C0(n403), .Y(
        Inst_forkAE_REG_TK2_0_N39) );
  AOI222XL U553 ( .A0(Inst_forkAE_KEY_INVERSE[37]), .A1(n193), .B0(n151), .B1(
        n208), .C0(n196), .C1(n404), .Y(n403) );
  XNOR2X1 U554 ( .A(n405), .B(randd[37]), .Y(n208) );
  CLKNAND2X2 U555 ( .A(IDtReg[37]), .B(MuxSel2), .Y(n405) );
  MXI2X1 U556 ( .A(n393), .B(n394), .S0(n406), .Y(n402) );
  NOR2BX1 U557 ( .AN(n210), .B(n407), .Y(n394) );
  AND2X1 U558 ( .A(n210), .B(n407), .Y(n393) );
  XOR2X1 U559 ( .A(n260), .B(n249), .Y(n407) );
  CLKINVX1 U560 ( .A(Inst_forkAE_KEY_INVERSE[3]), .Y(n249) );
  CLKINVX1 U561 ( .A(Inst_forkAE_KEY_INVERSE[2]), .Y(n260) );
  OAI221X1 U562 ( .A0(n233), .A1(n255), .B0(n142), .B1(n408), .C0(n409), .Y(
        Inst_forkAE_REG_TK2_0_N38) );
  AOI222XL U563 ( .A0(n196), .A1(n410), .B0(n210), .B1(n411), .C0(n154), .C1(
        n412), .Y(n409) );
  CLKINVX1 U564 ( .A(n253), .Y(n412) );
  XOR2X1 U565 ( .A(n413), .B(randd[36]), .Y(n253) );
  CLKNAND2X2 U566 ( .A(IDtReg[36]), .B(MuxSel2), .Y(n413) );
  XOR2X1 U567 ( .A(Inst_forkAE_KEY_INVERSE[2]), .B(n406), .Y(n411) );
  XOR2X1 U568 ( .A(Inst_forkAE_CURRENT_KEY_59_), .B(Inst_forkAE_KEY_INVERSE[1]), .Y(n406) );
  CLKINVX1 U569 ( .A(Inst_forkAE_KEY_INVERSE[13]), .Y(n408) );
  CLKINVX1 U570 ( .A(Inst_forkAE_KEY_INVERSE[36]), .Y(n255) );
  OAI2B11X1 U571 ( .A1N(Inst_forkAE_CURRENT_KEY_35_), .A0(n139), .B0(n414), 
        .C0(n415), .Y(Inst_forkAE_REG_TK2_0_N37) );
  AOI222XL U572 ( .A0(Inst_forkAE_KEY_INVERSE[35]), .A1(n193), .B0(n196), .B1(
        n416), .C0(n155), .C1(n330), .Y(n415) );
  XNOR2X1 U573 ( .A(n417), .B(randd[35]), .Y(n330) );
  CLKNAND2X2 U574 ( .A(IDtReg[35]), .B(MuxSel2), .Y(n417) );
  XOR2X1 U575 ( .A(n418), .B(n419), .Y(n416) );
  MXI2X1 U576 ( .A(n420), .B(n421), .S0(Inst_forkAE_CURRENT_KEY_47_), .Y(n414)
         );
  OAI211XL U577 ( .A0(n143), .A1(n355), .B0(n422), .C0(n423), .Y(
        Inst_forkAE_REG_TK2_0_N36) );
  AOI222XL U578 ( .A0(Inst_forkAE_KEY_INVERSE[34]), .A1(n193), .B0(n152), .B1(
        n400), .C0(n196), .C1(n418), .Y(n423) );
  XNOR2X1 U579 ( .A(n424), .B(randd[34]), .Y(n400) );
  CLKNAND2X2 U580 ( .A(IDtReg[34]), .B(MuxSel2), .Y(n424) );
  MXI2X1 U581 ( .A(n420), .B(n421), .S0(Inst_forkAE_KEY_INVERSE[21]), .Y(n422)
         );
  OAI211XL U582 ( .A0(n143), .A1(n354), .B0(n425), .C0(n426), .Y(
        Inst_forkAE_REG_TK2_0_N35) );
  AOI222XL U583 ( .A0(Inst_forkAE_KEY_INVERSE[33]), .A1(n193), .B0(n151), .B1(
        n427), .C0(n196), .C1(n428), .Y(n426) );
  MXI2X1 U584 ( .A(n420), .B(n421), .S0(n429), .Y(n425) );
  NOR2BX1 U585 ( .AN(n210), .B(n430), .Y(n421) );
  AND2X1 U586 ( .A(n210), .B(n430), .Y(n420) );
  XOR2X1 U587 ( .A(n347), .B(n343), .Y(n430) );
  CLKINVX1 U588 ( .A(Inst_forkAE_KEY_INVERSE[23]), .Y(n343) );
  CLKINVX1 U589 ( .A(Inst_forkAE_KEY_INVERSE[22]), .Y(n347) );
  OAI221X1 U590 ( .A0(n233), .A1(n431), .B0(n142), .B1(n432), .C0(n433), .Y(
        Inst_forkAE_REG_TK2_0_N34) );
  AOI222XL U591 ( .A0(n196), .A1(n434), .B0(n210), .B1(n435), .C0(n154), .C1(
        n436), .Y(n433) );
  CLKINVX1 U592 ( .A(n437), .Y(n436) );
  XOR2X1 U593 ( .A(Inst_forkAE_KEY_INVERSE[22]), .B(n429), .Y(n435) );
  XOR2X1 U594 ( .A(Inst_forkAE_CURRENT_KEY_47_), .B(
        Inst_forkAE_KEY_INVERSE[21]), .Y(n429) );
  CLKINVX1 U595 ( .A(Inst_forkAE_KEY_INVERSE[17]), .Y(n432) );
  OAI2B11X1 U596 ( .A1N(Inst_forkAE_KEY_INVERSE[63]), .A0(n139), .B0(n438), 
        .C0(n439), .Y(Inst_forkAE_REG_TK2_0_N33) );
  AOI222XL U597 ( .A0(Inst_forkAE_KEY_INVERSE[31]), .A1(n193), .B0(n151), .B1(
        n280), .C0(n196), .C1(n215), .Y(n439) );
  XNOR2X1 U598 ( .A(n440), .B(randd[63]), .Y(n215) );
  CLKNAND2X2 U599 ( .A(IDtReg[63]), .B(MuxSel2), .Y(n440) );
  XNOR2X1 U600 ( .A(n441), .B(randd[31]), .Y(n280) );
  CLKNAND2X2 U601 ( .A(IDtReg[31]), .B(MuxSel2), .Y(n441) );
  MXI2X1 U602 ( .A(n442), .B(n443), .S0(Inst_forkAE_KEY_INVERSE[43]), .Y(n438)
         );
  OAI2B11X1 U603 ( .A1N(Inst_forkAE_KEY_INVERSE[62]), .A0(n139), .B0(n444), 
        .C0(n445), .Y(Inst_forkAE_REG_TK2_0_N32) );
  AOI222XL U604 ( .A0(Inst_forkAE_KEY_INVERSE[30]), .A1(n193), .B0(n150), .B1(
        n291), .C0(n196), .C1(n223), .Y(n445) );
  XNOR2X1 U605 ( .A(n446), .B(randd[62]), .Y(n223) );
  CLKNAND2X2 U606 ( .A(IDtReg[62]), .B(MuxSel2), .Y(n446) );
  XNOR2X1 U607 ( .A(n447), .B(randd[30]), .Y(n291) );
  CLKNAND2X2 U608 ( .A(IDtReg[30]), .B(MuxSel2), .Y(n447) );
  MXI2X1 U609 ( .A(n442), .B(n443), .S0(Inst_forkAE_KEY_INVERSE[40]), .Y(n444)
         );
  OAI211XL U610 ( .A0(n143), .A1(n448), .B0(n449), .C0(n450), .Y(
        Inst_forkAE_REG_TK2_0_N31) );
  AOI222XL U611 ( .A0(Inst_forkAE_KEY_INVERSE[29]), .A1(n193), .B0(n152), .B1(
        n299), .C0(n196), .C1(n227), .Y(n450) );
  XNOR2X1 U612 ( .A(n451), .B(randd[61]), .Y(n227) );
  CLKNAND2X2 U613 ( .A(IDtReg[61]), .B(MuxSel2), .Y(n451) );
  XNOR2X1 U614 ( .A(n452), .B(randd[29]), .Y(n299) );
  CLKNAND2X2 U615 ( .A(IDtReg[29]), .B(MuxSel2), .Y(n452) );
  MXI2X1 U616 ( .A(n442), .B(n443), .S0(n453), .Y(n449) );
  NOR2BX1 U617 ( .AN(n210), .B(n454), .Y(n443) );
  AND2X1 U618 ( .A(n210), .B(n454), .Y(n442) );
  OAI221X1 U619 ( .A0(n240), .A1(n254), .B0(n141), .B1(n234), .C0(n455), .Y(
        Inst_forkAE_REG_TK2_0_N30) );
  AOI222XL U620 ( .A0(n153), .A1(n281), .B0(n193), .B1(n456), .C0(n210), .C1(
        n457), .Y(n455) );
  XOR2X1 U621 ( .A(Inst_forkAE_KEY_INVERSE[41]), .B(n453), .Y(n457) );
  XOR2X1 U622 ( .A(Inst_forkAE_KEY_INVERSE[43]), .B(
        Inst_forkAE_KEY_INVERSE[40]), .Y(n453) );
  XOR2X1 U623 ( .A(Inst_forkAE_KEY_INVERSE[31]), .B(
        Inst_forkAE_CURRENT_KEY_55_), .Y(n456) );
  XNOR2X1 U624 ( .A(n458), .B(randd[28]), .Y(n281) );
  CLKNAND2X2 U625 ( .A(IDtReg[28]), .B(MuxSel2), .Y(n458) );
  CLKINVX1 U626 ( .A(Inst_forkAE_KEY_INVERSE[60]), .Y(n234) );
  XOR2X1 U627 ( .A(n459), .B(randd[60]), .Y(n240) );
  CLKNAND2X2 U628 ( .A(IDtReg[60]), .B(MuxSel2), .Y(n459) );
  OAI211XL U629 ( .A0(n143), .A1(n460), .B0(n461), .C0(n462), .Y(
        Inst_forkAE_REG_TK2_0_N3) );
  AOI222XL U630 ( .A0(Inst_forkAE_KEY_INVERSE[1]), .A1(n193), .B0(n152), .B1(
        n272), .C0(n196), .C1(n427), .Y(n462) );
  XNOR2X1 U631 ( .A(n463), .B(randd[33]), .Y(n427) );
  CLKNAND2X2 U632 ( .A(IDtReg[33]), .B(MuxSel2), .Y(n463) );
  XNOR2X1 U633 ( .A(n464), .B(randd[1]), .Y(n272) );
  CLKNAND2X2 U634 ( .A(IDtReg[1]), .B(MuxSel2), .Y(n464) );
  MXI2X1 U635 ( .A(n332), .B(n333), .S0(n465), .Y(n461) );
  NOR2BX1 U636 ( .AN(n210), .B(n466), .Y(n333) );
  AND2X1 U637 ( .A(n210), .B(n466), .Y(n332) );
  OAI211XL U638 ( .A0(n143), .A1(n467), .B0(n468), .C0(n469), .Y(
        Inst_forkAE_REG_TK2_0_N29) );
  AOI222XL U639 ( .A0(Inst_forkAE_KEY_INVERSE[27]), .A1(n193), .B0(n151), .B1(
        n216), .C0(n196), .C1(n244), .Y(n469) );
  XNOR2X1 U640 ( .A(n470), .B(randd[59]), .Y(n244) );
  CLKNAND2X2 U641 ( .A(IDtReg[59]), .B(MuxSel2), .Y(n470) );
  XNOR2X1 U642 ( .A(n471), .B(randd[27]), .Y(n216) );
  CLKNAND2X2 U643 ( .A(IDtReg[27]), .B(MuxSel2), .Y(n471) );
  MXI2X1 U644 ( .A(n472), .B(n473), .S0(Inst_forkAE_KEY_INVERSE[39]), .Y(n468)
         );
  CLKINVX1 U645 ( .A(Inst_forkAE_KEY_INVERSE[59]), .Y(n467) );
  OAI211XL U646 ( .A0(n143), .A1(n474), .B0(n475), .C0(n476), .Y(
        Inst_forkAE_REG_TK2_0_N28) );
  AOI222XL U647 ( .A0(Inst_forkAE_KEY_INVERSE[26]), .A1(n193), .B0(n152), .B1(
        n228), .C0(n196), .C1(n252), .Y(n476) );
  XNOR2X1 U648 ( .A(n477), .B(randd[58]), .Y(n252) );
  CLKNAND2X2 U649 ( .A(IDtReg[58]), .B(MuxSel2), .Y(n477) );
  XNOR2X1 U650 ( .A(n478), .B(randd[26]), .Y(n228) );
  CLKNAND2X2 U651 ( .A(IDtReg[26]), .B(MuxSel2), .Y(n478) );
  MXI2X1 U652 ( .A(n472), .B(n473), .S0(Inst_forkAE_KEY_INVERSE[36]), .Y(n475)
         );
  OAI211XL U653 ( .A0(n143), .A1(n479), .B0(n480), .C0(n481), .Y(
        Inst_forkAE_REG_TK2_0_N27) );
  AOI222XL U654 ( .A0(Inst_forkAE_KEY_INVERSE[25]), .A1(n193), .B0(n152), .B1(
        n237), .C0(n196), .C1(n263), .Y(n481) );
  XNOR2X1 U655 ( .A(n482), .B(randd[57]), .Y(n263) );
  CLKNAND2X2 U656 ( .A(IDtReg[57]), .B(MuxSel2), .Y(n482) );
  XNOR2X1 U657 ( .A(n483), .B(randd[25]), .Y(n237) );
  CLKNAND2X2 U658 ( .A(IDtReg[25]), .B(MuxSel2), .Y(n483) );
  MXI2X1 U659 ( .A(n472), .B(n473), .S0(n484), .Y(n480) );
  NOR2BX1 U660 ( .AN(n210), .B(n485), .Y(n473) );
  AND2X1 U661 ( .A(n210), .B(n485), .Y(n472) );
  OAI221X1 U662 ( .A0(n275), .A1(n254), .B0(n142), .B1(n269), .C0(n486), .Y(
        Inst_forkAE_REG_TK2_0_N26) );
  AOI222XL U663 ( .A0(n153), .A1(n217), .B0(n193), .B1(n487), .C0(n210), .C1(
        n488), .Y(n486) );
  XOR2X1 U664 ( .A(Inst_forkAE_KEY_INVERSE[37]), .B(n484), .Y(n488) );
  XOR2X1 U665 ( .A(Inst_forkAE_KEY_INVERSE[39]), .B(
        Inst_forkAE_KEY_INVERSE[36]), .Y(n484) );
  XOR2X1 U666 ( .A(Inst_forkAE_KEY_INVERSE[27]), .B(
        Inst_forkAE_CURRENT_KEY_63_), .Y(n487) );
  XNOR2X1 U667 ( .A(n489), .B(randd[24]), .Y(n217) );
  CLKNAND2X2 U668 ( .A(IDtReg[24]), .B(MuxSel2), .Y(n489) );
  CLKINVX1 U669 ( .A(Inst_forkAE_KEY_INVERSE[56]), .Y(n269) );
  XOR2X1 U670 ( .A(n490), .B(randd[56]), .Y(n275) );
  CLKNAND2X2 U671 ( .A(IDtReg[56]), .B(MuxSel2), .Y(n490) );
  OAI2B11X1 U672 ( .A1N(Inst_forkAE_KEY_INVERSE[55]), .A0(n138), .B0(n491), 
        .C0(n492), .Y(Inst_forkAE_REG_TK2_0_N25) );
  AOI222XL U673 ( .A0(Inst_forkAE_KEY_INVERSE[23]), .A1(n193), .B0(n152), .B1(
        n339), .C0(n196), .C1(n279), .Y(n492) );
  XNOR2X1 U674 ( .A(n493), .B(randd[55]), .Y(n279) );
  CLKNAND2X2 U675 ( .A(IDtReg[55]), .B(MuxSel2), .Y(n493) );
  XNOR2X1 U676 ( .A(n494), .B(randd[23]), .Y(n339) );
  CLKNAND2X2 U677 ( .A(IDtReg[23]), .B(MuxSel2), .Y(n494) );
  MXI2X1 U678 ( .A(n495), .B(n496), .S0(Inst_forkAE_KEY_INVERSE[51]), .Y(n491)
         );
  OAI2B11X1 U679 ( .A1N(Inst_forkAE_KEY_INVERSE[54]), .A0(n139), .B0(n497), 
        .C0(n498), .Y(Inst_forkAE_REG_TK2_0_N24) );
  AOI222XL U680 ( .A0(Inst_forkAE_KEY_INVERSE[22]), .A1(n193), .B0(n151), .B1(
        n351), .C0(n196), .C1(n287), .Y(n498) );
  XNOR2X1 U681 ( .A(n499), .B(randd[54]), .Y(n287) );
  CLKNAND2X2 U682 ( .A(IDtReg[54]), .B(MuxSel2), .Y(n499) );
  XNOR2X1 U683 ( .A(n500), .B(randd[22]), .Y(n351) );
  CLKNAND2X2 U684 ( .A(IDtReg[22]), .B(MuxSel2), .Y(n500) );
  MXI2X1 U685 ( .A(n495), .B(n496), .S0(Inst_forkAE_KEY_INVERSE[48]), .Y(n497)
         );
  OAI211XL U686 ( .A0(n144), .A1(n501), .B0(n502), .C0(n503), .Y(
        Inst_forkAE_REG_TK2_0_N23) );
  AOI222XL U687 ( .A0(Inst_forkAE_KEY_INVERSE[21]), .A1(n193), .B0(n152), .B1(
        n359), .C0(n196), .C1(n290), .Y(n503) );
  XNOR2X1 U688 ( .A(n504), .B(randd[53]), .Y(n290) );
  CLKNAND2X2 U689 ( .A(IDtReg[53]), .B(MuxSel2), .Y(n504) );
  XNOR2X1 U690 ( .A(n505), .B(randd[21]), .Y(n359) );
  CLKNAND2X2 U691 ( .A(IDtReg[21]), .B(MuxSel2), .Y(n505) );
  MXI2X1 U692 ( .A(n495), .B(n496), .S0(n506), .Y(n502) );
  NOR2BX1 U693 ( .AN(n210), .B(n507), .Y(n496) );
  AND2X1 U694 ( .A(n210), .B(n507), .Y(n495) );
  OAI221X1 U695 ( .A0(n302), .A1(n254), .B0(n142), .B1(n296), .C0(n508), .Y(
        Inst_forkAE_REG_TK2_0_N22) );
  AOI222XL U696 ( .A0(n153), .A1(n340), .B0(n193), .B1(n509), .C0(n210), .C1(
        n510), .Y(n508) );
  XOR2X1 U697 ( .A(Inst_forkAE_KEY_INVERSE[49]), .B(n506), .Y(n510) );
  XOR2X1 U698 ( .A(Inst_forkAE_KEY_INVERSE[51]), .B(
        Inst_forkAE_KEY_INVERSE[48]), .Y(n506) );
  XOR2X1 U699 ( .A(Inst_forkAE_KEY_INVERSE[23]), .B(
        Inst_forkAE_CURRENT_KEY_47_), .Y(n509) );
  XNOR2X1 U700 ( .A(n511), .B(randd[20]), .Y(n340) );
  CLKNAND2X2 U701 ( .A(IDtReg[20]), .B(MuxSel2), .Y(n511) );
  CLKINVX1 U702 ( .A(Inst_forkAE_KEY_INVERSE[52]), .Y(n296) );
  XOR2X1 U703 ( .A(n512), .B(randd[52]), .Y(n302) );
  CLKNAND2X2 U704 ( .A(IDtReg[52]), .B(MuxSel2), .Y(n512) );
  OAI211XL U705 ( .A0(n144), .A1(n513), .B0(n514), .C0(n515), .Y(
        Inst_forkAE_REG_TK2_0_N21) );
  AOI222XL U706 ( .A0(Inst_forkAE_KEY_INVERSE[19]), .A1(n193), .B0(n152), .B1(
        n418), .C0(n196), .C1(n307), .Y(n515) );
  XNOR2X1 U707 ( .A(n516), .B(randd[51]), .Y(n307) );
  CLKNAND2X2 U708 ( .A(IDtReg[51]), .B(MuxSel2), .Y(n516) );
  XNOR2X1 U709 ( .A(n517), .B(randd[19]), .Y(n418) );
  CLKNAND2X2 U710 ( .A(IDtReg[19]), .B(MuxSel2), .Y(n517) );
  MXI2X1 U711 ( .A(n518), .B(n519), .S0(Inst_forkAE_KEY_INVERSE[55]), .Y(n514)
         );
  CLKINVX1 U712 ( .A(Inst_forkAE_KEY_INVERSE[51]), .Y(n513) );
  OAI211XL U713 ( .A0(n144), .A1(n520), .B0(n521), .C0(n522), .Y(
        Inst_forkAE_REG_TK2_0_N20) );
  AOI222XL U714 ( .A0(Inst_forkAE_KEY_INVERSE[18]), .A1(n193), .B0(n152), .B1(
        n428), .C0(n196), .C1(n314), .Y(n522) );
  XNOR2X1 U715 ( .A(n523), .B(randd[50]), .Y(n314) );
  CLKNAND2X2 U716 ( .A(IDtReg[50]), .B(MuxSel2), .Y(n523) );
  XNOR2X1 U717 ( .A(n524), .B(randd[18]), .Y(n428) );
  CLKNAND2X2 U718 ( .A(IDtReg[18]), .B(MuxSel2), .Y(n524) );
  MXI2X1 U719 ( .A(n518), .B(n519), .S0(Inst_forkAE_KEY_INVERSE[52]), .Y(n521)
         );
  OAI221X1 U720 ( .A0(n437), .A1(n254), .B0(n142), .B1(n431), .C0(n525), .Y(
        Inst_forkAE_REG_TK2_0_N2) );
  AOI222XL U721 ( .A0(n153), .A1(n246), .B0(n193), .B1(n526), .C0(n210), .C1(
        n527), .Y(n525) );
  XOR2X1 U722 ( .A(Inst_forkAE_KEY_INVERSE[45]), .B(n465), .Y(n527) );
  XOR2X1 U723 ( .A(Inst_forkAE_KEY_INVERSE[47]), .B(
        Inst_forkAE_KEY_INVERSE[44]), .Y(n465) );
  XOR2X1 U724 ( .A(Inst_forkAE_KEY_INVERSE[3]), .B(Inst_forkAE_CURRENT_KEY_59_), .Y(n526) );
  XNOR2X1 U725 ( .A(n528), .B(randd[0]), .Y(n246) );
  CLKNAND2X2 U726 ( .A(IDtReg[0]), .B(MuxSel2), .Y(n528) );
  XOR2X1 U727 ( .A(n529), .B(randd[32]), .Y(n437) );
  CLKNAND2X2 U728 ( .A(IDtReg[32]), .B(MuxSel2), .Y(n529) );
  OAI211XL U729 ( .A0(n144), .A1(n530), .B0(n531), .C0(n532), .Y(
        Inst_forkAE_REG_TK2_0_N19) );
  AOI222XL U730 ( .A0(Inst_forkAE_KEY_INVERSE[17]), .A1(n193), .B0(n153), .B1(
        n434), .C0(n196), .C1(n317), .Y(n532) );
  XNOR2X1 U731 ( .A(n533), .B(randd[49]), .Y(n317) );
  CLKNAND2X2 U732 ( .A(IDtReg[49]), .B(MuxSel2), .Y(n533) );
  XNOR2X1 U733 ( .A(n534), .B(randd[17]), .Y(n434) );
  CLKNAND2X2 U734 ( .A(IDtReg[17]), .B(MuxSel2), .Y(n534) );
  MXI2X1 U735 ( .A(n518), .B(n519), .S0(n535), .Y(n531) );
  NOR2BX1 U736 ( .AN(n210), .B(n536), .Y(n519) );
  AND2X1 U737 ( .A(n210), .B(n536), .Y(n518) );
  OAI221X1 U738 ( .A0(n327), .A1(n254), .B0(n142), .B1(n321), .C0(n537), .Y(
        Inst_forkAE_REG_TK2_0_N18) );
  AOI222XL U739 ( .A0(n153), .A1(n419), .B0(n193), .B1(n538), .C0(n210), .C1(
        n539), .Y(n537) );
  XOR2X1 U740 ( .A(Inst_forkAE_KEY_INVERSE[53]), .B(n535), .Y(n539) );
  XOR2X1 U741 ( .A(Inst_forkAE_KEY_INVERSE[55]), .B(
        Inst_forkAE_KEY_INVERSE[52]), .Y(n535) );
  XOR2X1 U742 ( .A(Inst_forkAE_KEY_INVERSE[19]), .B(
        Inst_forkAE_CURRENT_KEY_35_), .Y(n538) );
  XNOR2X1 U743 ( .A(n540), .B(randd[16]), .Y(n419) );
  CLKNAND2X2 U744 ( .A(IDtReg[16]), .B(MuxSel2), .Y(n540) );
  CLKINVX1 U745 ( .A(Inst_forkAE_KEY_INVERSE[48]), .Y(n321) );
  XOR2X1 U746 ( .A(n541), .B(randd[48]), .Y(n327) );
  CLKNAND2X2 U747 ( .A(IDtReg[48]), .B(MuxSel2), .Y(n541) );
  OAI211XL U748 ( .A0(n144), .A1(n542), .B0(n543), .C0(n544), .Y(
        Inst_forkAE_REG_TK2_0_N17) );
  AOI222XL U749 ( .A0(Inst_forkAE_KEY_INVERSE[15]), .A1(n193), .B0(n153), .B1(
        n391), .C0(n196), .C1(n338), .Y(n544) );
  XNOR2X1 U750 ( .A(n545), .B(randd[47]), .Y(n338) );
  CLKNAND2X2 U751 ( .A(IDtReg[47]), .B(MuxSel2), .Y(n545) );
  XNOR2X1 U752 ( .A(n546), .B(randd[15]), .Y(n391) );
  CLKNAND2X2 U753 ( .A(IDtReg[15]), .B(MuxSel2), .Y(n546) );
  MXI2X1 U754 ( .A(n547), .B(n548), .S0(Inst_forkAE_KEY_INVERSE[35]), .Y(n543)
         );
  CLKINVX1 U755 ( .A(Inst_forkAE_KEY_INVERSE[47]), .Y(n542) );
  OAI211XL U756 ( .A0(n144), .A1(n549), .B0(n550), .C0(n551), .Y(
        Inst_forkAE_REG_TK2_0_N16) );
  AOI222XL U757 ( .A0(Inst_forkAE_KEY_INVERSE[14]), .A1(n193), .B0(n152), .B1(
        n404), .C0(n196), .C1(n346), .Y(n551) );
  XNOR2X1 U758 ( .A(n552), .B(randd[46]), .Y(n346) );
  CLKNAND2X2 U759 ( .A(IDtReg[46]), .B(MuxSel2), .Y(n552) );
  XNOR2X1 U760 ( .A(n553), .B(randd[14]), .Y(n404) );
  CLKNAND2X2 U761 ( .A(IDtReg[14]), .B(MuxSel2), .Y(n553) );
  MXI2X1 U762 ( .A(n547), .B(n548), .S0(Inst_forkAE_KEY_INVERSE[32]), .Y(n550)
         );
  OAI211XL U763 ( .A0(n144), .A1(n554), .B0(n555), .C0(n556), .Y(
        Inst_forkAE_REG_TK2_0_N15) );
  AOI222XL U764 ( .A0(Inst_forkAE_KEY_INVERSE[13]), .A1(n193), .B0(n152), .B1(
        n410), .C0(n196), .C1(n350), .Y(n556) );
  XNOR2X1 U765 ( .A(n557), .B(randd[45]), .Y(n350) );
  CLKNAND2X2 U766 ( .A(IDtReg[45]), .B(MuxSel2), .Y(n557) );
  XNOR2X1 U767 ( .A(n558), .B(randd[13]), .Y(n410) );
  CLKNAND2X2 U768 ( .A(IDtReg[13]), .B(MuxSel2), .Y(n558) );
  MXI2X1 U769 ( .A(n547), .B(n548), .S0(n559), .Y(n555) );
  NOR2BX1 U770 ( .AN(n210), .B(n560), .Y(n548) );
  CLKINVX1 U771 ( .A(n561), .Y(n560) );
  NOR2BX1 U772 ( .AN(n210), .B(n561), .Y(n547) );
  OAI221X1 U773 ( .A0(n362), .A1(n254), .B0(n141), .B1(n356), .C0(n562), .Y(
        Inst_forkAE_REG_TK2_0_N14) );
  AOI222XL U774 ( .A0(n153), .A1(n392), .B0(n193), .B1(n563), .C0(n210), .C1(
        n564), .Y(n562) );
  XOR2X1 U775 ( .A(Inst_forkAE_KEY_INVERSE[33]), .B(n559), .Y(n564) );
  XOR2X1 U776 ( .A(Inst_forkAE_KEY_INVERSE[35]), .B(
        Inst_forkAE_KEY_INVERSE[32]), .Y(n559) );
  XOR2X1 U777 ( .A(Inst_forkAE_KEY_INVERSE[15]), .B(
        Inst_forkAE_CURRENT_KEY_39_), .Y(n563) );
  XNOR2X1 U778 ( .A(n565), .B(randd[12]), .Y(n392) );
  CLKNAND2X2 U779 ( .A(IDtReg[12]), .B(MuxSel2), .Y(n565) );
  CLKINVX1 U780 ( .A(Inst_forkAE_KEY_INVERSE[44]), .Y(n356) );
  XOR2X1 U781 ( .A(n566), .B(randd[44]), .Y(n362) );
  CLKNAND2X2 U782 ( .A(IDtReg[44]), .B(MuxSel2), .Y(n566) );
  OAI2B11X1 U783 ( .A1N(Inst_forkAE_KEY_INVERSE[43]), .A0(n139), .B0(n567), 
        .C0(n568), .Y(Inst_forkAE_REG_TK2_0_N13) );
  AOI222XL U784 ( .A0(Inst_forkAE_KEY_INVERSE[11]), .A1(n193), .B0(n153), .B1(
        n308), .C0(n196), .C1(n366), .Y(n568) );
  XNOR2X1 U785 ( .A(n569), .B(randd[43]), .Y(n366) );
  CLKNAND2X2 U786 ( .A(IDtReg[43]), .B(MuxSel2), .Y(n569) );
  XNOR2X1 U787 ( .A(n570), .B(randd[11]), .Y(n308) );
  CLKNAND2X2 U788 ( .A(IDtReg[11]), .B(MuxSel2), .Y(n570) );
  MXI2X1 U789 ( .A(n571), .B(n572), .S0(Inst_forkAE_KEY_INVERSE[63]), .Y(n567)
         );
  OAI211XL U790 ( .A0(n144), .A1(n573), .B0(n574), .C0(n575), .Y(
        Inst_forkAE_REG_TK2_0_N12) );
  AOI222XL U791 ( .A0(Inst_forkAE_KEY_INVERSE[10]), .A1(n193), .B0(n150), .B1(
        n318), .C0(n196), .C1(n372), .Y(n575) );
  XNOR2X1 U792 ( .A(n576), .B(randd[42]), .Y(n372) );
  CLKNAND2X2 U793 ( .A(IDtReg[42]), .B(MuxSel2), .Y(n576) );
  XNOR2X1 U794 ( .A(n577), .B(randd[10]), .Y(n318) );
  CLKNAND2X2 U795 ( .A(IDtReg[10]), .B(MuxSel2), .Y(n577) );
  MXI2X1 U796 ( .A(n571), .B(n572), .S0(Inst_forkAE_KEY_INVERSE[60]), .Y(n574)
         );
  OAI211XL U797 ( .A0(n144), .A1(n578), .B0(n579), .C0(n580), .Y(
        Inst_forkAE_REG_TK2_0_N11) );
  AOI222XL U798 ( .A0(Inst_forkAE_KEY_INVERSE[9]), .A1(n193), .B0(n153), .B1(
        n324), .C0(n196), .C1(n376), .Y(n580) );
  XNOR2X1 U799 ( .A(n581), .B(randd[41]), .Y(n376) );
  CLKNAND2X2 U800 ( .A(IDtReg[41]), .B(MuxSel2), .Y(n581) );
  XNOR2X1 U801 ( .A(n582), .B(randd[9]), .Y(n324) );
  CLKNAND2X2 U802 ( .A(IDtReg[9]), .B(MuxSel2), .Y(n582) );
  MXI2X1 U803 ( .A(n571), .B(n572), .S0(n583), .Y(n579) );
  NOR2BX1 U804 ( .AN(n210), .B(n584), .Y(n572) );
  AND2X1 U805 ( .A(n210), .B(n584), .Y(n571) );
  OAI221X1 U806 ( .A0(n385), .A1(n254), .B0(n142), .B1(n380), .C0(n585), .Y(
        Inst_forkAE_REG_TK2_0_N10) );
  AOI222XL U807 ( .A0(n153), .A1(n309), .B0(n193), .B1(n586), .C0(n210), .C1(
        n587), .Y(n585) );
  XOR2X1 U808 ( .A(Inst_forkAE_KEY_INVERSE[61]), .B(n583), .Y(n587) );
  XOR2X1 U809 ( .A(Inst_forkAE_KEY_INVERSE[63]), .B(
        Inst_forkAE_KEY_INVERSE[60]), .Y(n583) );
  XOR2X1 U810 ( .A(Inst_forkAE_KEY_INVERSE[11]), .B(
        Inst_forkAE_CURRENT_KEY_51_), .Y(n586) );
  XNOR2X1 U811 ( .A(n588), .B(randd[8]), .Y(n309) );
  CLKNAND2X2 U812 ( .A(IDtReg[8]), .B(MuxSel2), .Y(n588) );
  CLKINVX1 U813 ( .A(Inst_forkAE_KEY_INVERSE[40]), .Y(n380) );
  XOR2X1 U814 ( .A(n589), .B(randd[40]), .Y(n385) );
  CLKNAND2X2 U815 ( .A(IDtReg[40]), .B(MuxSel2), .Y(n589) );
  OAI2B11X1 U816 ( .A1N(Inst_forkAE_KEY_INVERSE[103]), .A0(n138), .B0(n590), 
        .C0(n591), .Y(Inst_forkAE_REG_TK2_N9) );
  AOI222XL U817 ( .A0(n592), .A1(n196), .B0(n193), .B1(n593), .C0(n594), .C1(
        n155), .Y(n591) );
  MXI2X1 U818 ( .A(n595), .B(n596), .S0(Inst_forkAE_KEY_INVERSE[122]), .Y(n590) );
  OAI2B11X1 U819 ( .A1N(Inst_forkAE_KEY_INVERSE[102]), .A0(n138), .B0(n597), 
        .C0(n598), .Y(Inst_forkAE_REG_TK2_N8) );
  AOI222XL U820 ( .A0(Inst_forkAE_KEY_INVERSE[70]), .A1(n193), .B0(n599), .B1(
        n158), .C0(n600), .C1(n196), .Y(n598) );
  MXI2X1 U821 ( .A(n595), .B(n596), .S0(Inst_forkAE_KEY_INVERSE[120]), .Y(n597) );
  OAI221X1 U822 ( .A0(n233), .A1(n601), .B0(n142), .B1(n602), .C0(n603), .Y(
        Inst_forkAE_REG_TK2_N7) );
  AOI222XL U823 ( .A0(n604), .A1(n196), .B0(n210), .B1(n605), .C0(n606), .C1(
        n155), .Y(n603) );
  XOR2X1 U824 ( .A(Inst_forkAE_KEY_INVERSE[122]), .B(n607), .Y(n605) );
  OAI2B11X1 U825 ( .A1N(Inst_forkAE_KEY_INVERSE[90]), .A0(n138), .B0(n608), 
        .C0(n609), .Y(Inst_forkAE_REG_TK2_N65) );
  AOI222XL U826 ( .A0(Inst_forkAE_KEY_INVERSE[127]), .A1(n193), .B0(n610), 
        .B1(n158), .C0(n611), .C1(n196), .Y(n609) );
  MXI2X1 U827 ( .A(n612), .B(n613), .S0(Inst_forkAE_KEY_INVERSE[69]), .Y(n608)
         );
  OAI211XL U828 ( .A0(n144), .A1(n614), .B0(n615), .C0(n616), .Y(
        Inst_forkAE_REG_TK2_N64) );
  AOI222XL U829 ( .A0(Inst_forkAE_KEY_INVERSE[126]), .A1(n193), .B0(n617), 
        .B1(n158), .C0(n618), .C1(n196), .Y(n616) );
  MXI2X1 U830 ( .A(n612), .B(n613), .S0(Inst_forkAE_CURRENT_KEY_104_), .Y(n615) );
  OAI221X1 U831 ( .A0(n233), .A1(n619), .B0(n141), .B1(n620), .C0(n621), .Y(
        Inst_forkAE_REG_TK2_N63) );
  AOI222XL U832 ( .A0(n622), .A1(n196), .B0(n210), .B1(n623), .C0(n624), .C1(
        n155), .Y(n621) );
  XOR2X1 U833 ( .A(Inst_forkAE_KEY_INVERSE[69]), .B(n593), .Y(n623) );
  XOR2X1 U834 ( .A(Inst_forkAE_CURRENT_KEY_104_), .B(
        Inst_forkAE_KEY_INVERSE[70]), .Y(n593) );
  OAI2B11X1 U835 ( .A1N(Inst_forkAE_CURRENT_KEY_124_), .A0(n138), .B0(n625), 
        .C0(n626), .Y(Inst_forkAE_REG_TK2_N62) );
  AOI222XL U836 ( .A0(Inst_forkAE_KEY_INVERSE[124]), .A1(n193), .B0(n196), 
        .B1(n627), .C0(n628), .C1(n155), .Y(n626) );
  XOR2X1 U837 ( .A(n611), .B(n629), .Y(n627) );
  MXI2X1 U838 ( .A(n612), .B(n613), .S0(Inst_forkAE_KEY_INVERSE[70]), .Y(n625)
         );
  NOR2BX1 U839 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[68]), .Y(n613) );
  NOR2BX1 U840 ( .AN(n210), .B(n630), .Y(n612) );
  OAI211XL U841 ( .A0(n144), .A1(n631), .B0(n632), .C0(n633), .Y(
        Inst_forkAE_REG_TK2_N61) );
  AOI222XL U842 ( .A0(Inst_forkAE_KEY_INVERSE[123]), .A1(n193), .B0(n634), 
        .B1(n158), .C0(n635), .C1(n196), .Y(n633) );
  MXI2X1 U843 ( .A(n636), .B(n637), .S0(Inst_forkAE_KEY_INVERSE[77]), .Y(n632)
         );
  OAI211XL U844 ( .A0(n144), .A1(n638), .B0(n639), .C0(n640), .Y(
        Inst_forkAE_REG_TK2_N60) );
  AOI222XL U845 ( .A0(Inst_forkAE_KEY_INVERSE[122]), .A1(n193), .B0(n641), 
        .B1(n158), .C0(n642), .C1(n196), .Y(n640) );
  MXI2X1 U846 ( .A(n636), .B(n637), .S0(Inst_forkAE_CURRENT_KEY_100_), .Y(n639) );
  OAI2B11X1 U847 ( .A1N(Inst_forkAE_KEY_INVERSE[100]), .A0(n137), .B0(n643), 
        .C0(n644), .Y(Inst_forkAE_REG_TK2_N6) );
  AOI222XL U848 ( .A0(Inst_forkAE_KEY_INVERSE[68]), .A1(n193), .B0(n645), .B1(
        n159), .C0(n646), .C1(n196), .Y(n644) );
  MXI2X1 U849 ( .A(n595), .B(n596), .S0(Inst_forkAE_KEY_INVERSE[123]), .Y(n643) );
  NOR2BX1 U850 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[121]), .Y(n596) );
  NOR2BX1 U851 ( .AN(n210), .B(n647), .Y(n595) );
  OAI221X1 U852 ( .A0(n233), .A1(n647), .B0(n141), .B1(n648), .C0(n649), .Y(
        Inst_forkAE_REG_TK2_N59) );
  AOI222XL U853 ( .A0(n650), .A1(n196), .B0(n210), .B1(n651), .C0(n652), .C1(
        n156), .Y(n649) );
  XOR2X1 U854 ( .A(Inst_forkAE_KEY_INVERSE[77]), .B(n653), .Y(n651) );
  OAI2B11X1 U855 ( .A1N(Inst_forkAE_CURRENT_KEY_120_), .A0(n138), .B0(n654), 
        .C0(n655), .Y(Inst_forkAE_REG_TK2_N58) );
  AOI222XL U856 ( .A0(Inst_forkAE_KEY_INVERSE[120]), .A1(n193), .B0(n196), 
        .B1(n656), .C0(n657), .C1(n155), .Y(n655) );
  XOR2X1 U857 ( .A(n635), .B(n658), .Y(n656) );
  MXI2X1 U858 ( .A(n636), .B(n637), .S0(Inst_forkAE_KEY_INVERSE[78]), .Y(n654)
         );
  NOR2BX1 U859 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[76]), .Y(n637) );
  NOR2BX1 U860 ( .AN(n210), .B(n659), .Y(n636) );
  OAI211XL U861 ( .A0(n144), .A1(n660), .B0(n661), .C0(n662), .Y(
        Inst_forkAE_REG_TK2_N57) );
  AOI222XL U862 ( .A0(Inst_forkAE_KEY_INVERSE[119]), .A1(n193), .B0(n663), 
        .B1(n158), .C0(n664), .C1(n196), .Y(n662) );
  MXI2X1 U863 ( .A(n665), .B(n666), .S0(Inst_forkAE_KEY_INVERSE[73]), .Y(n661)
         );
  OAI211XL U864 ( .A0(n144), .A1(n667), .B0(n668), .C0(n669), .Y(
        Inst_forkAE_REG_TK2_N56) );
  AOI222XL U865 ( .A0(Inst_forkAE_KEY_INVERSE[118]), .A1(n193), .B0(n670), 
        .B1(n158), .C0(n671), .C1(n196), .Y(n669) );
  MXI2X1 U866 ( .A(n665), .B(n666), .S0(Inst_forkAE_CURRENT_KEY_112_), .Y(n668) );
  OAI221X1 U867 ( .A0(n233), .A1(n672), .B0(n141), .B1(n673), .C0(n674), .Y(
        Inst_forkAE_REG_TK2_N55) );
  AOI222XL U868 ( .A0(n675), .A1(n196), .B0(n210), .B1(n676), .C0(n677), .C1(
        n155), .Y(n674) );
  XOR2X1 U869 ( .A(Inst_forkAE_KEY_INVERSE[73]), .B(n678), .Y(n676) );
  OAI2B11X1 U870 ( .A1N(Inst_forkAE_CURRENT_KEY_116_), .A0(n138), .B0(n679), 
        .C0(n680), .Y(Inst_forkAE_REG_TK2_N54) );
  AOI222XL U871 ( .A0(Inst_forkAE_KEY_INVERSE[116]), .A1(n193), .B0(n196), 
        .B1(n681), .C0(n682), .C1(n156), .Y(n680) );
  XOR2X1 U872 ( .A(n664), .B(n683), .Y(n681) );
  MXI2X1 U873 ( .A(n665), .B(n666), .S0(Inst_forkAE_KEY_INVERSE[74]), .Y(n679)
         );
  NOR2BX1 U874 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[72]), .Y(n666) );
  NOR2BX1 U875 ( .AN(n210), .B(n684), .Y(n665) );
  OAI2B11X1 U876 ( .A1N(Inst_forkAE_KEY_INVERSE[74]), .A0(n137), .B0(n685), 
        .C0(n686), .Y(Inst_forkAE_REG_TK2_N53) );
  AOI222XL U877 ( .A0(Inst_forkAE_KEY_INVERSE[115]), .A1(n193), .B0(n687), 
        .B1(n158), .C0(n688), .C1(n196), .Y(n686) );
  MXI2X1 U878 ( .A(n689), .B(n690), .S0(Inst_forkAE_KEY_INVERSE[93]), .Y(n685)
         );
  OAI211XL U879 ( .A0(n144), .A1(n691), .B0(n692), .C0(n693), .Y(
        Inst_forkAE_REG_TK2_N52) );
  AOI222XL U880 ( .A0(Inst_forkAE_KEY_INVERSE[114]), .A1(n193), .B0(n694), 
        .B1(n158), .C0(n695), .C1(n196), .Y(n693) );
  MXI2X1 U881 ( .A(n689), .B(n690), .S0(Inst_forkAE_CURRENT_KEY_116_), .Y(n692) );
  OAI221X1 U882 ( .A0(n233), .A1(n696), .B0(n141), .B1(n684), .C0(n697), .Y(
        Inst_forkAE_REG_TK2_N51) );
  AOI222XL U883 ( .A0(n698), .A1(n196), .B0(n210), .B1(n699), .C0(n700), .C1(
        n156), .Y(n697) );
  XOR2X1 U884 ( .A(Inst_forkAE_KEY_INVERSE[93]), .B(n701), .Y(n699) );
  CLKINVX1 U885 ( .A(Inst_forkAE_KEY_INVERSE[72]), .Y(n684) );
  OAI211XL U886 ( .A0(n144), .A1(n702), .B0(n703), .C0(n704), .Y(
        Inst_forkAE_REG_TK2_N50) );
  AOI222XL U887 ( .A0(Inst_forkAE_KEY_INVERSE[112]), .A1(n193), .B0(n196), 
        .B1(n705), .C0(n706), .C1(n155), .Y(n704) );
  XOR2X1 U888 ( .A(n688), .B(n707), .Y(n705) );
  MXI2X1 U889 ( .A(n689), .B(n690), .S0(Inst_forkAE_KEY_INVERSE[94]), .Y(n703)
         );
  NOR2BX1 U890 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[92]), .Y(n690) );
  NOR2BX1 U891 ( .AN(n210), .B(n673), .Y(n689) );
  CLKINVX1 U892 ( .A(Inst_forkAE_CURRENT_KEY_112_), .Y(n702) );
  OAI221X1 U893 ( .A0(n254), .A1(n708), .B0(n141), .B1(n709), .C0(n710), .Y(
        Inst_forkAE_REG_TK2_N5) );
  AOI222XL U894 ( .A0(n658), .A1(n154), .B0(n193), .B1(n711), .C0(n210), .C1(
        n712), .Y(n710) );
  XOR2X1 U895 ( .A(n713), .B(rand_in[3]), .Y(n658) );
  MX2X1 U896 ( .A(IDstReg[3]), .B(IDtReg[3]), .S0(DtSel), .Y(n713) );
  CLKINVX1 U897 ( .A(n714), .Y(n708) );
  OAI2B11X1 U898 ( .A1N(Inst_forkAE_KEY_INVERSE[86]), .A0(n138), .B0(n715), 
        .C0(n716), .Y(Inst_forkAE_REG_TK2_N49) );
  AOI222XL U899 ( .A0(Inst_forkAE_KEY_INVERSE[111]), .A1(n193), .B0(n717), 
        .B1(n158), .C0(n718), .C1(n196), .Y(n716) );
  MXI2X1 U900 ( .A(n719), .B(n720), .S0(Inst_forkAE_KEY_INVERSE[81]), .Y(n715)
         );
  OAI211XL U901 ( .A0(n144), .A1(n721), .B0(n722), .C0(n723), .Y(
        Inst_forkAE_REG_TK2_N48) );
  AOI222XL U902 ( .A0(Inst_forkAE_KEY_INVERSE[110]), .A1(n193), .B0(n724), 
        .B1(n158), .C0(n725), .C1(n196), .Y(n723) );
  MXI2X1 U903 ( .A(n719), .B(n720), .S0(Inst_forkAE_CURRENT_KEY_96_), .Y(n722)
         );
  OAI221X1 U904 ( .A0(n233), .A1(n726), .B0(n141), .B1(n727), .C0(n728), .Y(
        Inst_forkAE_REG_TK2_N47) );
  AOI222XL U905 ( .A0(n729), .A1(n196), .B0(n210), .B1(n730), .C0(n731), .C1(
        n156), .Y(n728) );
  XOR2X1 U906 ( .A(Inst_forkAE_KEY_INVERSE[81]), .B(n732), .Y(n730) );
  OAI2B11X1 U907 ( .A1N(Inst_forkAE_CURRENT_KEY_108_), .A0(n138), .B0(n733), 
        .C0(n734), .Y(Inst_forkAE_REG_TK2_N46) );
  AOI222XL U908 ( .A0(Inst_forkAE_KEY_INVERSE[108]), .A1(n193), .B0(n196), 
        .B1(n735), .C0(n736), .C1(n156), .Y(n734) );
  XOR2X1 U909 ( .A(n718), .B(n737), .Y(n735) );
  MXI2X1 U910 ( .A(n719), .B(n720), .S0(Inst_forkAE_KEY_INVERSE[82]), .Y(n733)
         );
  NOR2BX1 U911 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[80]), .Y(n720) );
  NOR2BX1 U912 ( .AN(n210), .B(n738), .Y(n719) );
  OAI211XL U913 ( .A0(n145), .A1(n739), .B0(n740), .C0(n741), .Y(
        Inst_forkAE_REG_TK2_N45) );
  AOI222XL U914 ( .A0(Inst_forkAE_KEY_INVERSE[107]), .A1(n193), .B0(n742), 
        .B1(n159), .C0(n599), .C1(n196), .Y(n741) );
  MXI2X1 U915 ( .A(n743), .B(n744), .S0(Inst_forkAE_KEY_INVERSE[89]), .Y(n740)
         );
  CLKINVX1 U916 ( .A(Inst_forkAE_KEY_INVERSE[70]), .Y(n739) );
  OAI211XL U917 ( .A0(n145), .A1(n601), .B0(n745), .C0(n746), .Y(
        Inst_forkAE_REG_TK2_N44) );
  AOI222XL U918 ( .A0(Inst_forkAE_KEY_INVERSE[106]), .A1(n193), .B0(n747), 
        .B1(n159), .C0(n606), .C1(n196), .Y(n746) );
  XOR2X1 U919 ( .A(n748), .B(rand_in[5]), .Y(n606) );
  MX2X1 U920 ( .A(IDstReg[5]), .B(IDtReg[5]), .S0(DtSel), .Y(n748) );
  MXI2X1 U921 ( .A(n743), .B(n744), .S0(Inst_forkAE_CURRENT_KEY_124_), .Y(n745) );
  OAI221X1 U922 ( .A0(n233), .A1(n749), .B0(n140), .B1(n630), .C0(n750), .Y(
        Inst_forkAE_REG_TK2_N43) );
  AOI222XL U923 ( .A0(n645), .A1(n196), .B0(n210), .B1(n751), .C0(n752), .C1(
        n157), .Y(n750) );
  XOR2X1 U924 ( .A(Inst_forkAE_KEY_INVERSE[89]), .B(n753), .Y(n751) );
  XOR2X1 U925 ( .A(n754), .B(rand_in[4]), .Y(n645) );
  MX2X1 U926 ( .A(IDstReg[4]), .B(IDtReg[4]), .S0(DtSel), .Y(n754) );
  CLKINVX1 U927 ( .A(Inst_forkAE_KEY_INVERSE[68]), .Y(n630) );
  OAI211XL U928 ( .A0(n145), .A1(n755), .B0(n756), .C0(n757), .Y(
        Inst_forkAE_REG_TK2_N42) );
  AOI222XL U929 ( .A0(Inst_forkAE_KEY_INVERSE[104]), .A1(n193), .B0(n196), 
        .B1(n758), .C0(n759), .C1(n156), .Y(n757) );
  XOR2X1 U930 ( .A(n594), .B(n599), .Y(n758) );
  XOR2X1 U931 ( .A(n760), .B(rand_in[6]), .Y(n599) );
  MX2X1 U932 ( .A(IDstReg[6]), .B(IDtReg[6]), .S0(DtSel), .Y(n760) );
  XOR2X1 U933 ( .A(n761), .B(rand_in[7]), .Y(n594) );
  MX2X1 U934 ( .A(IDstReg[7]), .B(IDtReg[7]), .S0(DtSel), .Y(n761) );
  MXI2X1 U935 ( .A(n743), .B(n744), .S0(Inst_forkAE_KEY_INVERSE[90]), .Y(n756)
         );
  NOR2BX1 U936 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[88]), .Y(n744) );
  NOR2BX1 U937 ( .AN(n210), .B(n620), .Y(n743) );
  CLKINVX1 U938 ( .A(Inst_forkAE_KEY_INVERSE[88]), .Y(n620) );
  CLKINVX1 U939 ( .A(Inst_forkAE_CURRENT_KEY_104_), .Y(n755) );
  OAI211XL U940 ( .A0(n145), .A1(n762), .B0(n763), .C0(n764), .Y(
        Inst_forkAE_REG_TK2_N41) );
  AOI222XL U941 ( .A0(Inst_forkAE_KEY_INVERSE[103]), .A1(n193), .B0(n592), 
        .B1(n158), .C0(n765), .C1(n196), .Y(n764) );
  XOR2X1 U942 ( .A(n766), .B(rand_in[39]), .Y(n592) );
  MX2X1 U943 ( .A(IDstReg[39]), .B(IDtReg[39]), .S0(DtSel), .Y(n766) );
  MXI2X1 U944 ( .A(n767), .B(n768), .S0(Inst_forkAE_KEY_INVERSE[65]), .Y(n763)
         );
  OAI211XL U945 ( .A0(n145), .A1(n769), .B0(n770), .C0(n771), .Y(
        Inst_forkAE_REG_TK2_N40) );
  AOI222XL U946 ( .A0(Inst_forkAE_KEY_INVERSE[102]), .A1(n193), .B0(n600), 
        .B1(n159), .C0(n772), .C1(n196), .Y(n771) );
  XOR2X1 U947 ( .A(n773), .B(rand_in[38]), .Y(n600) );
  MX2X1 U948 ( .A(IDstReg[38]), .B(IDtReg[38]), .S0(DtSel), .Y(n773) );
  MXI2X1 U949 ( .A(n767), .B(n768), .S0(Inst_forkAE_CURRENT_KEY_120_), .Y(n770) );
  OAI221X1 U950 ( .A0(n233), .A1(n631), .B0(n140), .B1(n774), .C0(n775), .Y(
        Inst_forkAE_REG_TK2_N4) );
  AOI222XL U951 ( .A0(n776), .A1(n196), .B0(n210), .B1(n777), .C0(n635), .C1(
        n155), .Y(n775) );
  XOR2X1 U952 ( .A(n778), .B(rand_in[2]), .Y(n635) );
  MX2X1 U953 ( .A(IDstReg[2]), .B(IDtReg[2]), .S0(DtSel), .Y(n778) );
  XOR2X1 U954 ( .A(Inst_forkAE_KEY_INVERSE[109]), .B(
        Inst_forkAE_KEY_INVERSE[108]), .Y(n777) );
  CLKINVX1 U955 ( .A(Inst_forkAE_KEY_INVERSE[98]), .Y(n774) );
  CLKINVX1 U956 ( .A(Inst_forkAE_KEY_INVERSE[66]), .Y(n631) );
  OAI221X1 U957 ( .A0(n233), .A1(n602), .B0(n140), .B1(n659), .C0(n779), .Y(
        Inst_forkAE_REG_TK2_N39) );
  AOI222XL U958 ( .A0(n780), .A1(n196), .B0(n210), .B1(n781), .C0(n604), .C1(
        n157), .Y(n779) );
  XOR2X1 U959 ( .A(n782), .B(rand_in[37]), .Y(n604) );
  MX2X1 U960 ( .A(IDstReg[37]), .B(IDtReg[37]), .S0(DtSel), .Y(n782) );
  XOR2X1 U961 ( .A(Inst_forkAE_KEY_INVERSE[65]), .B(n711), .Y(n781) );
  XOR2X1 U962 ( .A(Inst_forkAE_CURRENT_KEY_120_), .B(
        Inst_forkAE_KEY_INVERSE[66]), .Y(n711) );
  OAI211XL U963 ( .A0(n145), .A1(n783), .B0(n784), .C0(n785), .Y(
        Inst_forkAE_REG_TK2_N38) );
  AOI222XL U964 ( .A0(Inst_forkAE_KEY_INVERSE[100]), .A1(n193), .B0(n196), 
        .B1(n786), .C0(n646), .C1(n156), .Y(n785) );
  XOR2X1 U965 ( .A(n787), .B(rand_in[36]), .Y(n646) );
  MX2X1 U966 ( .A(IDstReg[36]), .B(IDtReg[36]), .S0(DtSel), .Y(n787) );
  XOR2X1 U967 ( .A(n765), .B(n788), .Y(n786) );
  MXI2X1 U968 ( .A(n767), .B(n768), .S0(Inst_forkAE_KEY_INVERSE[66]), .Y(n784)
         );
  NOR2BX1 U969 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[64]), .Y(n768) );
  NOR2BX1 U970 ( .AN(n210), .B(n648), .Y(n767) );
  CLKINVX1 U971 ( .A(Inst_forkAE_CURRENT_KEY_100_), .Y(n783) );
  OAI211XL U972 ( .A0(n145), .A1(n789), .B0(n790), .C0(n791), .Y(
        Inst_forkAE_REG_TK2_N37) );
  AOI222XL U973 ( .A0(Inst_forkAE_KEY_INVERSE[99]), .A1(n193), .B0(n714), .B1(
        n158), .C0(n792), .C1(n196), .Y(n791) );
  XOR2X1 U974 ( .A(n793), .B(rand_in[35]), .Y(n714) );
  MX2X1 U975 ( .A(IDstReg[35]), .B(IDtReg[35]), .S0(DtSel), .Y(n793) );
  MXI2X1 U976 ( .A(n794), .B(n795), .S0(Inst_forkAE_KEY_INVERSE[85]), .Y(n790)
         );
  CLKINVX1 U977 ( .A(Inst_forkAE_KEY_INVERSE[82]), .Y(n789) );
  OAI211XL U978 ( .A0(n145), .A1(n796), .B0(n797), .C0(n798), .Y(
        Inst_forkAE_REG_TK2_N36) );
  AOI222XL U979 ( .A0(Inst_forkAE_KEY_INVERSE[98]), .A1(n193), .B0(n776), .B1(
        n159), .C0(n799), .C1(n196), .Y(n798) );
  XOR2X1 U980 ( .A(n800), .B(rand_in[34]), .Y(n776) );
  MX2X1 U981 ( .A(IDstReg[34]), .B(IDtReg[34]), .S0(DtSel), .Y(n800) );
  MXI2X1 U982 ( .A(n794), .B(n795), .S0(Inst_forkAE_CURRENT_KEY_108_), .Y(n797) );
  OAI221X1 U983 ( .A0(n233), .A1(n801), .B0(n140), .B1(n738), .C0(n802), .Y(
        Inst_forkAE_REG_TK2_N35) );
  AOI222XL U984 ( .A0(n803), .A1(n196), .B0(n210), .B1(n804), .C0(n805), .C1(
        n156), .Y(n802) );
  XOR2X1 U985 ( .A(Inst_forkAE_KEY_INVERSE[85]), .B(n806), .Y(n804) );
  CLKINVX1 U986 ( .A(Inst_forkAE_KEY_INVERSE[80]), .Y(n738) );
  OAI211XL U987 ( .A0(n145), .A1(n807), .B0(n808), .C0(n809), .Y(
        Inst_forkAE_REG_TK2_N34) );
  AOI222XL U988 ( .A0(Inst_forkAE_KEY_INVERSE[96]), .A1(n193), .B0(n196), .B1(
        n810), .C0(n811), .C1(n156), .Y(n809) );
  XOR2X1 U989 ( .A(n792), .B(n812), .Y(n810) );
  MXI2X1 U990 ( .A(n794), .B(n795), .S0(Inst_forkAE_KEY_INVERSE[86]), .Y(n808)
         );
  NOR2BX1 U991 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[84]), .Y(n795) );
  NOR2BX1 U992 ( .AN(n210), .B(n727), .Y(n794) );
  CLKINVX1 U993 ( .A(Inst_forkAE_KEY_INVERSE[84]), .Y(n727) );
  CLKINVX1 U994 ( .A(Inst_forkAE_CURRENT_KEY_96_), .Y(n807) );
  OAI221X1 U995 ( .A0(n254), .A1(n813), .B0(n140), .B1(n814), .C0(n815), .Y(
        Inst_forkAE_REG_TK2_N33) );
  AOI222XL U996 ( .A0(n683), .A1(n154), .B0(n210), .B1(n816), .C0(n193), .C1(
        n701), .Y(n815) );
  XOR2X1 U997 ( .A(Inst_forkAE_CURRENT_KEY_116_), .B(
        Inst_forkAE_KEY_INVERSE[94]), .Y(n701) );
  XOR2X1 U998 ( .A(n817), .B(rand_in[31]), .Y(n683) );
  MX2X1 U999 ( .A(IDstReg[31]), .B(IDtReg[31]), .S0(DtSel), .Y(n817) );
  CLKINVX1 U1000 ( .A(Inst_forkAE_KEY_INVERSE[127]), .Y(n814) );
  CLKINVX1 U1001 ( .A(n610), .Y(n813) );
  XOR2X1 U1002 ( .A(n818), .B(rand_in[63]), .Y(n610) );
  MX2X1 U1003 ( .A(IDstReg[63]), .B(IDtReg[63]), .S0(DtSel), .Y(n818) );
  OAI221X1 U1004 ( .A0(n233), .A1(n660), .B0(n140), .B1(n819), .C0(n820), .Y(
        Inst_forkAE_REG_TK2_N32) );
  AOI222XL U1005 ( .A0(n617), .A1(n196), .B0(n210), .B1(n821), .C0(n664), .C1(
        n157), .Y(n820) );
  XOR2X1 U1006 ( .A(n822), .B(rand_in[30]), .Y(n664) );
  MX2X1 U1007 ( .A(IDstReg[30]), .B(IDtReg[30]), .S0(DtSel), .Y(n822) );
  XOR2X1 U1008 ( .A(Inst_forkAE_KEY_INVERSE[105]), .B(
        Inst_forkAE_KEY_INVERSE[104]), .Y(n821) );
  XOR2X1 U1009 ( .A(n823), .B(rand_in[62]), .Y(n617) );
  MX2X1 U1010 ( .A(IDstReg[62]), .B(IDtReg[62]), .S0(DtSel), .Y(n823) );
  CLKINVX1 U1011 ( .A(Inst_forkAE_KEY_INVERSE[126]), .Y(n819) );
  CLKINVX1 U1012 ( .A(Inst_forkAE_KEY_INVERSE[94]), .Y(n660) );
  OAI221X1 U1013 ( .A0(n233), .A1(n667), .B0(n140), .B1(n619), .C0(n824), .Y(
        Inst_forkAE_REG_TK2_N31) );
  AOI222XL U1014 ( .A0(n624), .A1(n196), .B0(n210), .B1(n825), .C0(n671), .C1(
        n156), .Y(n824) );
  XOR2X1 U1015 ( .A(n826), .B(rand_in[29]), .Y(n671) );
  MX2X1 U1016 ( .A(IDstReg[29]), .B(IDtReg[29]), .S0(DtSel), .Y(n826) );
  XOR2X1 U1017 ( .A(Inst_forkAE_KEY_INVERSE[106]), .B(n827), .Y(n825) );
  XOR2X1 U1018 ( .A(n828), .B(rand_in[61]), .Y(n624) );
  MX2X1 U1019 ( .A(IDstReg[61]), .B(IDtReg[61]), .S0(DtSel), .Y(n828) );
  CLKINVX1 U1020 ( .A(Inst_forkAE_KEY_INVERSE[93]), .Y(n667) );
  OAI221X1 U1021 ( .A0(n233), .A1(n673), .B0(n141), .B1(n829), .C0(n830), .Y(
        Inst_forkAE_REG_TK2_N30) );
  AOI222XL U1022 ( .A0(n628), .A1(n196), .B0(n210), .B1(n831), .C0(n675), .C1(
        n157), .Y(n830) );
  XOR2X1 U1023 ( .A(n832), .B(rand_in[28]), .Y(n675) );
  MX2X1 U1024 ( .A(IDstReg[28]), .B(IDtReg[28]), .S0(DtSel), .Y(n832) );
  XOR2X1 U1025 ( .A(Inst_forkAE_KEY_INVERSE[107]), .B(
        Inst_forkAE_KEY_INVERSE[105]), .Y(n831) );
  XOR2X1 U1026 ( .A(n833), .B(rand_in[60]), .Y(n628) );
  MX2X1 U1027 ( .A(IDstReg[60]), .B(IDtReg[60]), .S0(DtSel), .Y(n833) );
  CLKINVX1 U1028 ( .A(Inst_forkAE_KEY_INVERSE[92]), .Y(n673) );
  OAI221X1 U1029 ( .A0(n233), .A1(n638), .B0(n140), .B1(n801), .C0(n834), .Y(
        Inst_forkAE_REG_TK2_N3) );
  AOI222XL U1030 ( .A0(n805), .A1(n196), .B0(n210), .B1(n835), .C0(n642), .C1(
        n156), .Y(n834) );
  XOR2X1 U1031 ( .A(n836), .B(rand_in[1]), .Y(n642) );
  MX2X1 U1032 ( .A(IDstReg[1]), .B(IDtReg[1]), .S0(DtSel), .Y(n836) );
  XOR2X1 U1033 ( .A(Inst_forkAE_KEY_INVERSE[110]), .B(n837), .Y(n835) );
  XOR2X1 U1034 ( .A(n838), .B(rand_in[33]), .Y(n805) );
  MX2X1 U1035 ( .A(IDstReg[33]), .B(IDtReg[33]), .S0(DtSel), .Y(n838) );
  CLKINVX1 U1036 ( .A(Inst_forkAE_KEY_INVERSE[97]), .Y(n801) );
  CLKINVX1 U1037 ( .A(Inst_forkAE_KEY_INVERSE[65]), .Y(n638) );
  OAI211XL U1038 ( .A0(n145), .A1(n839), .B0(n840), .C0(n841), .Y(
        Inst_forkAE_REG_TK2_N29) );
  AOI222XL U1039 ( .A0(n634), .A1(n196), .B0(n193), .B1(n753), .C0(n629), .C1(
        n157), .Y(n841) );
  XOR2X1 U1040 ( .A(n842), .B(rand_in[27]), .Y(n629) );
  MX2X1 U1041 ( .A(IDstReg[27]), .B(IDtReg[27]), .S0(DtSel), .Y(n842) );
  XOR2X1 U1042 ( .A(Inst_forkAE_CURRENT_KEY_124_), .B(
        Inst_forkAE_KEY_INVERSE[90]), .Y(n753) );
  XOR2X1 U1043 ( .A(n843), .B(rand_in[59]), .Y(n634) );
  MX2X1 U1044 ( .A(IDstReg[59]), .B(IDtReg[59]), .S0(DtSel), .Y(n843) );
  MXI2X1 U1045 ( .A(n844), .B(n845), .S0(Inst_forkAE_KEY_INVERSE[102]), .Y(
        n840) );
  CLKINVX1 U1046 ( .A(Inst_forkAE_KEY_INVERSE[123]), .Y(n839) );
  OAI211XL U1047 ( .A0(n145), .A1(n846), .B0(n847), .C0(n848), .Y(
        Inst_forkAE_REG_TK2_N28) );
  AOI222XL U1048 ( .A0(Inst_forkAE_KEY_INVERSE[90]), .A1(n193), .B0(n611), 
        .B1(n159), .C0(n641), .C1(n196), .Y(n848) );
  XOR2X1 U1049 ( .A(n849), .B(rand_in[58]), .Y(n641) );
  MX2X1 U1050 ( .A(IDstReg[58]), .B(IDtReg[58]), .S0(DtSel), .Y(n849) );
  XOR2X1 U1051 ( .A(n850), .B(rand_in[26]), .Y(n611) );
  MX2X1 U1052 ( .A(IDstReg[26]), .B(IDtReg[26]), .S0(DtSel), .Y(n850) );
  MXI2X1 U1053 ( .A(n844), .B(n845), .S0(Inst_forkAE_KEY_INVERSE[100]), .Y(
        n847) );
  CLKINVX1 U1054 ( .A(Inst_forkAE_KEY_INVERSE[122]), .Y(n846) );
  OAI221X1 U1055 ( .A0(n233), .A1(n614), .B0(n140), .B1(n647), .C0(n851), .Y(
        Inst_forkAE_REG_TK2_N27) );
  AOI222XL U1056 ( .A0(n652), .A1(n196), .B0(n210), .B1(n852), .C0(n618), .C1(
        n157), .Y(n851) );
  XOR2X1 U1057 ( .A(n853), .B(rand_in[25]), .Y(n618) );
  MX2X1 U1058 ( .A(IDstReg[25]), .B(IDtReg[25]), .S0(DtSel), .Y(n853) );
  XOR2X1 U1059 ( .A(Inst_forkAE_KEY_INVERSE[102]), .B(n854), .Y(n852) );
  XOR2X1 U1060 ( .A(n855), .B(rand_in[57]), .Y(n652) );
  MX2X1 U1061 ( .A(IDstReg[57]), .B(IDtReg[57]), .S0(DtSel), .Y(n855) );
  CLKINVX1 U1062 ( .A(Inst_forkAE_KEY_INVERSE[89]), .Y(n614) );
  OAI2B11X1 U1063 ( .A1N(Inst_forkAE_KEY_INVERSE[120]), .A0(n137), .B0(n856), 
        .C0(n857), .Y(Inst_forkAE_REG_TK2_N26) );
  AOI222XL U1064 ( .A0(Inst_forkAE_KEY_INVERSE[88]), .A1(n193), .B0(n622), 
        .B1(n159), .C0(n657), .C1(n196), .Y(n857) );
  XOR2X1 U1065 ( .A(n858), .B(rand_in[56]), .Y(n657) );
  MX2X1 U1066 ( .A(IDstReg[56]), .B(IDtReg[56]), .S0(DtSel), .Y(n858) );
  XOR2X1 U1067 ( .A(n859), .B(rand_in[24]), .Y(n622) );
  MX2X1 U1068 ( .A(IDstReg[24]), .B(IDtReg[24]), .S0(DtSel), .Y(n859) );
  MXI2X1 U1069 ( .A(n844), .B(n845), .S0(Inst_forkAE_KEY_INVERSE[103]), .Y(
        n856) );
  NOR2BX1 U1070 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[101]), .Y(n845) );
  NOR2BX1 U1071 ( .AN(n210), .B(n602), .Y(n844) );
  OAI2B11X1 U1072 ( .A1N(Inst_forkAE_KEY_INVERSE[119]), .A0(n137), .B0(n860), 
        .C0(n861), .Y(Inst_forkAE_REG_TK2_N25) );
  AOI222XL U1073 ( .A0(n663), .A1(n196), .B0(n193), .B1(n806), .C0(n737), .C1(
        n157), .Y(n861) );
  XOR2X1 U1074 ( .A(n862), .B(rand_in[23]), .Y(n737) );
  MX2X1 U1075 ( .A(IDstReg[23]), .B(IDtReg[23]), .S0(DtSel), .Y(n862) );
  XOR2X1 U1076 ( .A(Inst_forkAE_CURRENT_KEY_108_), .B(
        Inst_forkAE_KEY_INVERSE[86]), .Y(n806) );
  XOR2X1 U1077 ( .A(n863), .B(rand_in[55]), .Y(n663) );
  MX2X1 U1078 ( .A(IDstReg[55]), .B(IDtReg[55]), .S0(DtSel), .Y(n863) );
  MXI2X1 U1079 ( .A(n864), .B(n865), .S0(Inst_forkAE_KEY_INVERSE[114]), .Y(
        n860) );
  OAI2B11X1 U1080 ( .A1N(Inst_forkAE_KEY_INVERSE[118]), .A0(n137), .B0(n866), 
        .C0(n867), .Y(Inst_forkAE_REG_TK2_N24) );
  AOI222XL U1081 ( .A0(Inst_forkAE_KEY_INVERSE[86]), .A1(n193), .B0(n718), 
        .B1(n159), .C0(n670), .C1(n196), .Y(n867) );
  XOR2X1 U1082 ( .A(n868), .B(rand_in[54]), .Y(n670) );
  MX2X1 U1083 ( .A(IDstReg[54]), .B(IDtReg[54]), .S0(DtSel), .Y(n868) );
  XOR2X1 U1084 ( .A(n869), .B(rand_in[22]), .Y(n718) );
  MX2X1 U1085 ( .A(IDstReg[22]), .B(IDtReg[22]), .S0(DtSel), .Y(n869) );
  MXI2X1 U1086 ( .A(n864), .B(n865), .S0(Inst_forkAE_KEY_INVERSE[112]), .Y(
        n866) );
  OAI221X1 U1087 ( .A0(n233), .A1(n721), .B0(n140), .B1(n672), .C0(n870), .Y(
        Inst_forkAE_REG_TK2_N23) );
  AOI222XL U1088 ( .A0(n677), .A1(n196), .B0(n210), .B1(n871), .C0(n725), .C1(
        n157), .Y(n870) );
  XOR2X1 U1089 ( .A(n872), .B(rand_in[21]), .Y(n725) );
  MX2X1 U1090 ( .A(IDstReg[21]), .B(IDtReg[21]), .S0(DtSel), .Y(n872) );
  XOR2X1 U1091 ( .A(Inst_forkAE_KEY_INVERSE[114]), .B(n873), .Y(n871) );
  XOR2X1 U1092 ( .A(n874), .B(rand_in[53]), .Y(n677) );
  MX2X1 U1093 ( .A(IDstReg[53]), .B(IDtReg[53]), .S0(DtSel), .Y(n874) );
  CLKINVX1 U1094 ( .A(Inst_forkAE_KEY_INVERSE[85]), .Y(n721) );
  OAI2B11X1 U1095 ( .A1N(Inst_forkAE_KEY_INVERSE[116]), .A0(n137), .B0(n875), 
        .C0(n876), .Y(Inst_forkAE_REG_TK2_N22) );
  AOI222XL U1096 ( .A0(Inst_forkAE_KEY_INVERSE[84]), .A1(n193), .B0(n729), 
        .B1(n159), .C0(n682), .C1(n196), .Y(n876) );
  XOR2X1 U1097 ( .A(n877), .B(rand_in[52]), .Y(n682) );
  MX2X1 U1098 ( .A(IDstReg[52]), .B(IDtReg[52]), .S0(DtSel), .Y(n877) );
  XOR2X1 U1099 ( .A(n878), .B(rand_in[20]), .Y(n729) );
  MX2X1 U1100 ( .A(IDstReg[20]), .B(IDtReg[20]), .S0(DtSel), .Y(n878) );
  MXI2X1 U1101 ( .A(n864), .B(n865), .S0(Inst_forkAE_KEY_INVERSE[115]), .Y(
        n875) );
  NOR2BX1 U1102 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[113]), .Y(n865) );
  NOR2BX1 U1103 ( .AN(n210), .B(n696), .Y(n864) );
  OAI211XL U1104 ( .A0(n145), .A1(n879), .B0(n880), .C0(n881), .Y(
        Inst_forkAE_REG_TK2_N21) );
  AOI222XL U1105 ( .A0(n687), .A1(n196), .B0(n193), .B1(n732), .C0(n812), .C1(
        n157), .Y(n881) );
  XOR2X1 U1106 ( .A(n882), .B(rand_in[19]), .Y(n812) );
  MX2X1 U1107 ( .A(IDstReg[19]), .B(IDtReg[19]), .S0(DtSel), .Y(n882) );
  XOR2X1 U1108 ( .A(Inst_forkAE_CURRENT_KEY_96_), .B(
        Inst_forkAE_KEY_INVERSE[82]), .Y(n732) );
  XOR2X1 U1109 ( .A(n883), .B(rand_in[51]), .Y(n687) );
  MX2X1 U1110 ( .A(IDstReg[51]), .B(IDtReg[51]), .S0(DtSel), .Y(n883) );
  MXI2X1 U1111 ( .A(n884), .B(n885), .S0(Inst_forkAE_KEY_INVERSE[118]), .Y(
        n880) );
  CLKINVX1 U1112 ( .A(Inst_forkAE_KEY_INVERSE[115]), .Y(n879) );
  OAI211XL U1113 ( .A0(n145), .A1(n886), .B0(n887), .C0(n888), .Y(
        Inst_forkAE_REG_TK2_N20) );
  AOI222XL U1114 ( .A0(Inst_forkAE_KEY_INVERSE[82]), .A1(n193), .B0(n792), 
        .B1(n159), .C0(n694), .C1(n196), .Y(n888) );
  XOR2X1 U1115 ( .A(n889), .B(rand_in[50]), .Y(n694) );
  MX2X1 U1116 ( .A(IDstReg[50]), .B(IDtReg[50]), .S0(DtSel), .Y(n889) );
  XOR2X1 U1117 ( .A(n890), .B(rand_in[18]), .Y(n792) );
  MX2X1 U1118 ( .A(IDstReg[18]), .B(IDtReg[18]), .S0(DtSel), .Y(n890) );
  MXI2X1 U1119 ( .A(n884), .B(n885), .S0(Inst_forkAE_KEY_INVERSE[116]), .Y(
        n887) );
  CLKINVX1 U1120 ( .A(Inst_forkAE_KEY_INVERSE[114]), .Y(n886) );
  OAI221X1 U1121 ( .A0(n233), .A1(n648), .B0(n139), .B1(n891), .C0(n892), .Y(
        Inst_forkAE_REG_TK2_N2) );
  AOI222XL U1122 ( .A0(n811), .A1(n196), .B0(n210), .B1(n893), .C0(n650), .C1(
        n157), .Y(n892) );
  XOR2X1 U1123 ( .A(n894), .B(rand_in[0]), .Y(n650) );
  MX2X1 U1124 ( .A(IDstReg[0]), .B(IDtReg[0]), .S0(DtSel), .Y(n894) );
  XOR2X1 U1125 ( .A(Inst_forkAE_KEY_INVERSE[111]), .B(
        Inst_forkAE_KEY_INVERSE[109]), .Y(n893) );
  XOR2X1 U1126 ( .A(n895), .B(rand_in[32]), .Y(n811) );
  MX2X1 U1127 ( .A(IDstReg[32]), .B(IDtReg[32]), .S0(DtSel), .Y(n895) );
  CLKINVX1 U1128 ( .A(Inst_forkAE_KEY_INVERSE[64]), .Y(n648) );
  OAI221X1 U1129 ( .A0(n233), .A1(n796), .B0(n139), .B1(n696), .C0(n896), .Y(
        Inst_forkAE_REG_TK2_N19) );
  AOI222XL U1130 ( .A0(n700), .A1(n196), .B0(n210), .B1(n897), .C0(n799), .C1(
        n156), .Y(n896) );
  XOR2X1 U1131 ( .A(n898), .B(rand_in[17]), .Y(n799) );
  MX2X1 U1132 ( .A(IDstReg[17]), .B(IDtReg[17]), .S0(DtSel), .Y(n898) );
  XOR2X1 U1133 ( .A(Inst_forkAE_KEY_INVERSE[118]), .B(n899), .Y(n897) );
  XOR2X1 U1134 ( .A(n900), .B(rand_in[49]), .Y(n700) );
  MX2X1 U1135 ( .A(IDstReg[49]), .B(IDtReg[49]), .S0(DtSel), .Y(n900) );
  CLKINVX1 U1136 ( .A(Inst_forkAE_KEY_INVERSE[81]), .Y(n796) );
  OAI2B11X1 U1137 ( .A1N(Inst_forkAE_KEY_INVERSE[112]), .A0(n137), .B0(n901), 
        .C0(n902), .Y(Inst_forkAE_REG_TK2_N18) );
  AOI222XL U1138 ( .A0(Inst_forkAE_KEY_INVERSE[80]), .A1(n193), .B0(n803), 
        .B1(n159), .C0(n706), .C1(n196), .Y(n902) );
  XOR2X1 U1139 ( .A(n903), .B(rand_in[48]), .Y(n706) );
  MX2X1 U1140 ( .A(IDstReg[48]), .B(IDtReg[48]), .S0(DtSel), .Y(n903) );
  XOR2X1 U1141 ( .A(n904), .B(rand_in[16]), .Y(n803) );
  MX2X1 U1142 ( .A(IDstReg[16]), .B(IDtReg[16]), .S0(DtSel), .Y(n904) );
  MXI2X1 U1143 ( .A(n884), .B(n885), .S0(Inst_forkAE_KEY_INVERSE[119]), .Y(
        n901) );
  NOR2BX1 U1144 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[117]), .Y(n885) );
  NOR2BX1 U1145 ( .AN(n210), .B(n672), .Y(n884) );
  OAI221X1 U1146 ( .A0(n254), .A1(n905), .B0(n139), .B1(n906), .C0(n907), .Y(
        Inst_forkAE_REG_TK2_N17) );
  AOI222XL U1147 ( .A0(n788), .A1(n153), .B0(n210), .B1(n908), .C0(n193), .C1(
        n653), .Y(n907) );
  XOR2X1 U1148 ( .A(Inst_forkAE_CURRENT_KEY_100_), .B(
        Inst_forkAE_KEY_INVERSE[78]), .Y(n653) );
  XOR2X1 U1149 ( .A(n909), .B(rand_in[15]), .Y(n788) );
  MX2X1 U1150 ( .A(IDstReg[15]), .B(IDtReg[15]), .S0(DtSel), .Y(n909) );
  CLKINVX1 U1151 ( .A(Inst_forkAE_KEY_INVERSE[111]), .Y(n906) );
  CLKINVX1 U1152 ( .A(n717), .Y(n905) );
  XOR2X1 U1153 ( .A(n910), .B(rand_in[47]), .Y(n717) );
  MX2X1 U1154 ( .A(IDstReg[47]), .B(IDtReg[47]), .S0(DtSel), .Y(n910) );
  CLKINVX1 U1155 ( .A(n196), .Y(n254) );
  OAI221X1 U1156 ( .A0(n233), .A1(n762), .B0(n141), .B1(n911), .C0(n912), .Y(
        Inst_forkAE_REG_TK2_N16) );
  AOI222XL U1157 ( .A0(n724), .A1(n196), .B0(n210), .B1(n913), .C0(n765), .C1(
        n157), .Y(n912) );
  XOR2X1 U1158 ( .A(n914), .B(rand_in[14]), .Y(n765) );
  MX2X1 U1159 ( .A(IDstReg[14]), .B(IDtReg[14]), .S0(DtSel), .Y(n914) );
  XOR2X1 U1160 ( .A(Inst_forkAE_KEY_INVERSE[97]), .B(
        Inst_forkAE_KEY_INVERSE[96]), .Y(n913) );
  XOR2X1 U1161 ( .A(n915), .B(rand_in[46]), .Y(n724) );
  MX2X1 U1162 ( .A(IDstReg[46]), .B(IDtReg[46]), .S0(DtSel), .Y(n915) );
  CLKINVX1 U1163 ( .A(Inst_forkAE_KEY_INVERSE[110]), .Y(n911) );
  CLKINVX1 U1164 ( .A(Inst_forkAE_KEY_INVERSE[78]), .Y(n762) );
  OAI221X1 U1165 ( .A0(n233), .A1(n769), .B0(n140), .B1(n726), .C0(n916), .Y(
        Inst_forkAE_REG_TK2_N15) );
  AOI222XL U1166 ( .A0(n731), .A1(n196), .B0(n210), .B1(n917), .C0(n772), .C1(
        n156), .Y(n916) );
  XOR2X1 U1167 ( .A(n918), .B(rand_in[13]), .Y(n772) );
  MX2X1 U1168 ( .A(IDstReg[13]), .B(IDtReg[13]), .S0(DtSel), .Y(n918) );
  XOR2X1 U1169 ( .A(Inst_forkAE_KEY_INVERSE[98]), .B(n919), .Y(n917) );
  XOR2X1 U1170 ( .A(n920), .B(rand_in[45]), .Y(n731) );
  MX2X1 U1171 ( .A(IDstReg[45]), .B(IDtReg[45]), .S0(DtSel), .Y(n920) );
  CLKINVX1 U1172 ( .A(Inst_forkAE_KEY_INVERSE[109]), .Y(n726) );
  CLKINVX1 U1173 ( .A(Inst_forkAE_KEY_INVERSE[77]), .Y(n769) );
  OAI221X1 U1174 ( .A0(n233), .A1(n659), .B0(n139), .B1(n921), .C0(n922), .Y(
        Inst_forkAE_REG_TK2_N14) );
  AOI222XL U1175 ( .A0(n736), .A1(n196), .B0(n210), .B1(n923), .C0(n780), .C1(
        n157), .Y(n922) );
  XOR2X1 U1176 ( .A(n924), .B(rand_in[12]), .Y(n780) );
  MX2X1 U1177 ( .A(IDstReg[12]), .B(IDtReg[12]), .S0(DtSel), .Y(n924) );
  XOR2X1 U1178 ( .A(Inst_forkAE_KEY_INVERSE[99]), .B(
        Inst_forkAE_KEY_INVERSE[97]), .Y(n923) );
  XOR2X1 U1179 ( .A(n925), .B(rand_in[44]), .Y(n736) );
  MX2X1 U1180 ( .A(IDstReg[44]), .B(IDtReg[44]), .S0(DtSel), .Y(n925) );
  CLKINVX1 U1181 ( .A(Inst_forkAE_KEY_INVERSE[108]), .Y(n921) );
  CLKINVX1 U1182 ( .A(Inst_forkAE_KEY_INVERSE[76]), .Y(n659) );
  OAI211XL U1183 ( .A0(n145), .A1(n926), .B0(n927), .C0(n928), .Y(
        Inst_forkAE_REG_TK2_N13) );
  AOI222XL U1184 ( .A0(n742), .A1(n196), .B0(n193), .B1(n678), .C0(n707), .C1(
        n157), .Y(n928) );
  XOR2X1 U1185 ( .A(n929), .B(rand_in[11]), .Y(n707) );
  MX2X1 U1186 ( .A(IDstReg[11]), .B(IDtReg[11]), .S0(DtSel), .Y(n929) );
  XOR2X1 U1187 ( .A(Inst_forkAE_CURRENT_KEY_112_), .B(
        Inst_forkAE_KEY_INVERSE[74]), .Y(n678) );
  XOR2X1 U1188 ( .A(n930), .B(rand_in[43]), .Y(n742) );
  MX2X1 U1189 ( .A(IDstReg[43]), .B(IDtReg[43]), .S0(DtSel), .Y(n930) );
  MXI2X1 U1190 ( .A(n931), .B(n932), .S0(Inst_forkAE_KEY_INVERSE[126]), .Y(
        n927) );
  CLKINVX1 U1191 ( .A(Inst_forkAE_KEY_INVERSE[107]), .Y(n926) );
  OAI2B11X1 U1192 ( .A1N(Inst_forkAE_KEY_INVERSE[106]), .A0(n137), .B0(n933), 
        .C0(n934), .Y(Inst_forkAE_REG_TK2_N12) );
  AOI222XL U1193 ( .A0(Inst_forkAE_KEY_INVERSE[74]), .A1(n193), .B0(n688), 
        .B1(n159), .C0(n747), .C1(n196), .Y(n934) );
  XOR2X1 U1194 ( .A(n935), .B(rand_in[42]), .Y(n747) );
  MX2X1 U1195 ( .A(IDstReg[42]), .B(IDtReg[42]), .S0(DtSel), .Y(n935) );
  XOR2X1 U1196 ( .A(n936), .B(rand_in[10]), .Y(n688) );
  MX2X1 U1197 ( .A(IDstReg[10]), .B(IDtReg[10]), .S0(DtSel), .Y(n936) );
  MXI2X1 U1198 ( .A(n931), .B(n932), .S0(Inst_forkAE_KEY_INVERSE[124]), .Y(
        n933) );
  OAI221X1 U1199 ( .A0(n233), .A1(n691), .B0(n139), .B1(n749), .C0(n937), .Y(
        Inst_forkAE_REG_TK2_N11) );
  AOI222XL U1200 ( .A0(n752), .A1(n196), .B0(n210), .B1(n938), .C0(n695), .C1(
        n158), .Y(n937) );
  XOR2X1 U1201 ( .A(n939), .B(rand_in[9]), .Y(n695) );
  MX2X1 U1202 ( .A(IDstReg[9]), .B(IDtReg[9]), .S0(DtSel), .Y(n939) );
  XOR2X1 U1203 ( .A(Inst_forkAE_KEY_INVERSE[126]), .B(n940), .Y(n938) );
  XOR2X1 U1204 ( .A(n941), .B(rand_in[41]), .Y(n752) );
  MX2X1 U1205 ( .A(IDstReg[41]), .B(IDtReg[41]), .S0(DtSel), .Y(n941) );
  CLKINVX1 U1206 ( .A(Inst_forkAE_KEY_INVERSE[105]), .Y(n749) );
  CLKINVX1 U1207 ( .A(Inst_forkAE_KEY_INVERSE[73]), .Y(n691) );
  OAI2B11X1 U1208 ( .A1N(Inst_forkAE_KEY_INVERSE[104]), .A0(n137), .B0(n942), 
        .C0(n943), .Y(Inst_forkAE_REG_TK2_N10) );
  AOI222XL U1209 ( .A0(Inst_forkAE_KEY_INVERSE[72]), .A1(n193), .B0(n698), 
        .B1(n159), .C0(n759), .C1(n196), .Y(n943) );
  XOR2X1 U1210 ( .A(n946), .B(rand_in[40]), .Y(n759) );
  MX2X1 U1211 ( .A(IDstReg[40]), .B(IDtReg[40]), .S0(DtSel), .Y(n946) );
  NOR2X1 U1212 ( .A(n944), .B(n947), .Y(n194) );
  XOR2X1 U1213 ( .A(n948), .B(rand_in[8]), .Y(n698) );
  MX2X1 U1214 ( .A(IDstReg[8]), .B(IDtReg[8]), .S0(DtSel), .Y(n948) );
  CLKINVX1 U1215 ( .A(n945), .Y(n947) );
  MXI2X1 U1216 ( .A(n931), .B(n932), .S0(Inst_forkAE_KEY_INVERSE[127]), .Y(
        n942) );
  NOR2BX1 U1217 ( .AN(n210), .B(Inst_forkAE_KEY_INVERSE[125]), .Y(n932) );
  NOR2BX1 U1218 ( .AN(n210), .B(n619), .Y(n931) );
  NAND3XL U1219 ( .A(n949), .B(n950), .C(n951), .Y(n945) );
  OAI21X1 U1220 ( .A0(n184), .A1(GO), .B0(n951), .Y(n944) );
  CLKNAND2X2 U1221 ( .A(n952), .B(n950), .Y(n190) );
  XOR2X1 U1222 ( .A(n953), .B(n954), .Y(n952) );
  XOR2X1 U1223 ( .A(Inst_forkAE_FSM_X_state_2_), .B(n955), .Y(n954) );
  OAI22X1 U1224 ( .A0(n956), .A1(n957), .B0(n955), .B1(n958), .Y(n953) );
  OA21X1 U1225 ( .A0(Inst_forkAE_FSM_X_state_1_), .A1(n957), .B0(n951), .Y(
        n955) );
  OAI221X1 U1226 ( .A0(C1[7]), .A1(n959), .B0(n960), .B1(n961), .C0(n962), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N9) );
  AOI22XL U1227 ( .A0(PLAINTEXT[7]), .A1(n963), .B0(n964), .B1(n965), .Y(n962)
         );
  CLKINVX1 U1228 ( .A(n966), .Y(n965) );
  OAI221X1 U1229 ( .A0(n959), .A1(n967), .B0(n968), .B1(n961), .C0(n969), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N8) );
  AOI22XL U1230 ( .A0(PLAINTEXT[6]), .A1(n963), .B0(n964), .B1(n970), .Y(n969)
         );
  CLKINVX1 U1231 ( .A(n971), .Y(n970) );
  OAI221X1 U1232 ( .A0(n959), .A1(n972), .B0(n973), .B1(n961), .C0(n974), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N7) );
  AOI22XL U1233 ( .A0(PLAINTEXT[5]), .A1(n963), .B0(n964), .B1(n975), .Y(n974)
         );
  OAI221X1 U1234 ( .A0(n959), .A1(n976), .B0(n961), .B1(n977), .C0(n978), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N65) );
  AOI22XL U1235 ( .A0(PLAINTEXT[63]), .A1(n963), .B0(n979), .B1(n964), .Y(n978) );
  OAI221X1 U1236 ( .A0(n959), .A1(n980), .B0(n981), .B1(n961), .C0(n982), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N64) );
  AOI22XL U1237 ( .A0(PLAINTEXT[62]), .A1(n963), .B0(n964), .B1(n983), .Y(n982) );
  CLKINVX1 U1238 ( .A(n984), .Y(n983) );
  CLKINVX1 U1239 ( .A(C1[62]), .Y(n980) );
  OAI221X1 U1240 ( .A0(n959), .A1(n985), .B0(n986), .B1(n961), .C0(n987), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N63) );
  AOI22XL U1241 ( .A0(PLAINTEXT[61]), .A1(n963), .B0(n964), .B1(n988), .Y(n987) );
  CLKINVX1 U1242 ( .A(n989), .Y(n988) );
  OAI221X1 U1243 ( .A0(C1[60]), .A1(n959), .B0(n990), .B1(n961), .C0(n991), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N62) );
  AOI22XL U1244 ( .A0(PLAINTEXT[60]), .A1(n963), .B0(n992), .B1(n964), .Y(n991) );
  OAI221X1 U1245 ( .A0(n959), .A1(n993), .B0(n994), .B1(n961), .C0(n995), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N61) );
  AOI22XL U1246 ( .A0(PLAINTEXT[59]), .A1(n963), .B0(n964), .B1(n996), .Y(n995) );
  CLKINVX1 U1247 ( .A(n997), .Y(n996) );
  CLKINVX1 U1248 ( .A(C1[59]), .Y(n993) );
  OAI221X1 U1249 ( .A0(n959), .A1(n998), .B0(n999), .B1(n961), .C0(n1000), .Y(
        Inst_forkAE_REG_INTERNAL_STATE_N60) );
  AOI22XL U1250 ( .A0(PLAINTEXT[58]), .A1(n963), .B0(n964), .B1(n1001), .Y(
        n1000) );
  CLKINVX1 U1251 ( .A(n1002), .Y(n1001) );
  CLKINVX1 U1252 ( .A(C1[58]), .Y(n998) );
  OAI221X1 U1253 ( .A0(n959), .A1(n1003), .B0(n1004), .B1(n961), .C0(n1005), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N6) );
  AOI22XL U1254 ( .A0(PLAINTEXT[4]), .A1(n963), .B0(n964), .B1(n1006), .Y(
        n1005) );
  CLKINVX1 U1255 ( .A(n1007), .Y(n1006) );
  OAI221X1 U1256 ( .A0(C1[57]), .A1(n959), .B0(n1008), .B1(n961), .C0(n1009), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N59) );
  AOI22XL U1257 ( .A0(PLAINTEXT[57]), .A1(n963), .B0(n964), .B1(n1010), .Y(
        n1009) );
  CLKINVX1 U1258 ( .A(n1011), .Y(n1010) );
  OAI221X1 U1259 ( .A0(n959), .A1(n1012), .B0(n1013), .B1(n961), .C0(n1014), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N58) );
  AOI22XL U1260 ( .A0(PLAINTEXT[56]), .A1(n963), .B0(n964), .B1(n1015), .Y(
        n1014) );
  CLKINVX1 U1261 ( .A(n1016), .Y(n1015) );
  CLKINVX1 U1262 ( .A(C1[56]), .Y(n1012) );
  OAI221X1 U1263 ( .A0(n959), .A1(n1017), .B0(n1018), .B1(n961), .C0(n1019), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N57) );
  AOI22XL U1264 ( .A0(PLAINTEXT[55]), .A1(n963), .B0(n964), .B1(n1020), .Y(
        n1019) );
  CLKINVX1 U1265 ( .A(n1021), .Y(n1020) );
  CLKINVX1 U1266 ( .A(C1[55]), .Y(n1017) );
  OAI221X1 U1267 ( .A0(C1[54]), .A1(n959), .B0(n1022), .B1(n961), .C0(n1023), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N56) );
  AOI22XL U1268 ( .A0(PLAINTEXT[54]), .A1(n963), .B0(n1024), .B1(n964), .Y(
        n1023) );
  OAI221X1 U1269 ( .A0(n959), .A1(n1025), .B0(n1026), .B1(n961), .C0(n1027), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N55) );
  AOI22XL U1270 ( .A0(PLAINTEXT[53]), .A1(n963), .B0(n964), .B1(n1028), .Y(
        n1027) );
  CLKINVX1 U1271 ( .A(n1029), .Y(n1028) );
  OAI221X1 U1272 ( .A0(n959), .A1(n1030), .B0(n1031), .B1(n961), .C0(n1032), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N54) );
  AOI22XL U1273 ( .A0(PLAINTEXT[52]), .A1(n963), .B0(n964), .B1(n1033), .Y(
        n1032) );
  CLKINVX1 U1274 ( .A(n1034), .Y(n1033) );
  CLKINVX1 U1275 ( .A(C1[52]), .Y(n1030) );
  OAI221X1 U1276 ( .A0(C1[51]), .A1(n959), .B0(n1035), .B1(n961), .C0(n1036), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N53) );
  AOI22XL U1277 ( .A0(PLAINTEXT[51]), .A1(n963), .B0(n964), .B1(n1037), .Y(
        n1036) );
  CLKINVX1 U1278 ( .A(n1038), .Y(n1037) );
  OAI221X1 U1279 ( .A0(n959), .A1(n1039), .B0(n1040), .B1(n961), .C0(n1041), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N52) );
  AOI22XL U1280 ( .A0(PLAINTEXT[50]), .A1(n963), .B0(n964), .B1(n1042), .Y(
        n1041) );
  CLKINVX1 U1281 ( .A(n1043), .Y(n1042) );
  CLKINVX1 U1282 ( .A(C1[50]), .Y(n1039) );
  OAI221X1 U1283 ( .A0(n959), .A1(n1044), .B0(n1045), .B1(n961), .C0(n1046), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N51) );
  AOI22XL U1284 ( .A0(PLAINTEXT[49]), .A1(n963), .B0(n964), .B1(n1047), .Y(
        n1046) );
  CLKINVX1 U1285 ( .A(n1048), .Y(n1047) );
  OAI221X1 U1286 ( .A0(C1[48]), .A1(n959), .B0(n1049), .B1(n961), .C0(n1050), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N50) );
  AOI22XL U1287 ( .A0(PLAINTEXT[48]), .A1(n963), .B0(n964), .B1(n1051), .Y(
        n1050) );
  CLKINVX1 U1288 ( .A(n1052), .Y(n1051) );
  OAI221X1 U1289 ( .A0(n959), .A1(n1053), .B0(n1054), .B1(n961), .C0(n1055), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N5) );
  AOI22XL U1290 ( .A0(PLAINTEXT[3]), .A1(n963), .B0(n964), .B1(n1056), .Y(
        n1055) );
  CLKINVX1 U1291 ( .A(n1057), .Y(n1056) );
  OAI221X1 U1292 ( .A0(n959), .A1(n1058), .B0(n961), .B1(n1059), .C0(n1060), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N49) );
  AOI22XL U1293 ( .A0(PLAINTEXT[47]), .A1(n963), .B0(n964), .B1(n1061), .Y(
        n1060) );
  CLKINVX1 U1294 ( .A(n1062), .Y(n1061) );
  CLKINVX1 U1295 ( .A(C1[47]), .Y(n1058) );
  OAI221X1 U1296 ( .A0(n959), .A1(n1063), .B0(n1064), .B1(n961), .C0(n1065), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N48) );
  AOI22XL U1297 ( .A0(PLAINTEXT[46]), .A1(n963), .B0(n1066), .B1(n964), .Y(
        n1065) );
  CLKINVX1 U1298 ( .A(C1[46]), .Y(n1063) );
  OAI221X1 U1299 ( .A0(C1[45]), .A1(n959), .B0(n1067), .B1(n961), .C0(n1068), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N47) );
  AOI22XL U1300 ( .A0(PLAINTEXT[45]), .A1(n963), .B0(n964), .B1(n1069), .Y(
        n1068) );
  CLKINVX1 U1301 ( .A(n1070), .Y(n1069) );
  OAI221X1 U1302 ( .A0(C1[44]), .A1(n959), .B0(n1071), .B1(n961), .C0(n1072), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N46) );
  AOI22XL U1303 ( .A0(PLAINTEXT[44]), .A1(n963), .B0(n964), .B1(n1073), .Y(
        n1072) );
  CLKINVX1 U1304 ( .A(n1074), .Y(n1073) );
  OAI221X1 U1305 ( .A0(n959), .A1(n1075), .B0(n1076), .B1(n961), .C0(n1077), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N45) );
  AOI22XL U1306 ( .A0(PLAINTEXT[43]), .A1(n963), .B0(n964), .B1(n1078), .Y(
        n1077) );
  CLKINVX1 U1307 ( .A(n1079), .Y(n1078) );
  CLKINVX1 U1308 ( .A(C1[43]), .Y(n1075) );
  OAI221X1 U1309 ( .A0(C1[42]), .A1(n959), .B0(n1080), .B1(n961), .C0(n1081), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N44) );
  AOI22XL U1310 ( .A0(PLAINTEXT[42]), .A1(n963), .B0(n964), .B1(n1082), .Y(
        n1081) );
  CLKINVX1 U1311 ( .A(n1083), .Y(n1082) );
  OAI221X1 U1312 ( .A0(C1[41]), .A1(n959), .B0(n1084), .B1(n961), .C0(n1085), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N43) );
  AOI22XL U1313 ( .A0(PLAINTEXT[41]), .A1(n963), .B0(n964), .B1(n1086), .Y(
        n1085) );
  CLKINVX1 U1314 ( .A(n1087), .Y(n1086) );
  OAI221X1 U1315 ( .A0(n959), .A1(n1088), .B0(n1089), .B1(n961), .C0(n1090), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N42) );
  AOI22XL U1316 ( .A0(PLAINTEXT[40]), .A1(n963), .B0(n964), .B1(n1091), .Y(
        n1090) );
  CLKINVX1 U1317 ( .A(n1092), .Y(n1091) );
  OAI221X1 U1318 ( .A0(C1[39]), .A1(n959), .B0(n1093), .B1(n961), .C0(n1094), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N41) );
  AOI22XL U1319 ( .A0(PLAINTEXT[39]), .A1(n963), .B0(n964), .B1(n1095), .Y(
        n1094) );
  CLKINVX1 U1320 ( .A(n1096), .Y(n1095) );
  OAI221X1 U1321 ( .A0(C1[38]), .A1(n959), .B0(n1097), .B1(n961), .C0(n1098), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N40) );
  AOI22XL U1322 ( .A0(PLAINTEXT[38]), .A1(n963), .B0(n964), .B1(n1099), .Y(
        n1098) );
  CLKINVX1 U1323 ( .A(n1100), .Y(n1099) );
  OAI221X1 U1324 ( .A0(n959), .A1(n1101), .B0(n1102), .B1(n961), .C0(n1103), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N4) );
  AOI22XL U1325 ( .A0(PLAINTEXT[2]), .A1(n963), .B0(n964), .B1(n1104), .Y(
        n1103) );
  CLKINVX1 U1326 ( .A(n1105), .Y(n1104) );
  OAI221X1 U1327 ( .A0(n959), .A1(n1106), .B0(n961), .B1(n1107), .C0(n1108), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N39) );
  AOI22XL U1328 ( .A0(PLAINTEXT[37]), .A1(n963), .B0(n964), .B1(n1109), .Y(
        n1108) );
  CLKINVX1 U1329 ( .A(n1110), .Y(n1109) );
  OAI221X1 U1330 ( .A0(C1[36]), .A1(n959), .B0(n1111), .B1(n961), .C0(n1112), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N38) );
  AOI22XL U1331 ( .A0(PLAINTEXT[36]), .A1(n963), .B0(n964), .B1(n1113), .Y(
        n1112) );
  CLKINVX1 U1332 ( .A(n1114), .Y(n1113) );
  OAI221X1 U1333 ( .A0(C1[35]), .A1(n959), .B0(n1115), .B1(n961), .C0(n1116), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N37) );
  AOI22XL U1334 ( .A0(PLAINTEXT[35]), .A1(n963), .B0(n964), .B1(n1117), .Y(
        n1116) );
  CLKINVX1 U1335 ( .A(n1118), .Y(n1117) );
  OAI221X1 U1336 ( .A0(n959), .A1(n1119), .B0(n1120), .B1(n961), .C0(n1121), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N36) );
  AOI22XL U1337 ( .A0(PLAINTEXT[34]), .A1(n963), .B0(n964), .B1(n1122), .Y(
        n1121) );
  CLKINVX1 U1338 ( .A(n1123), .Y(n1122) );
  OAI221X1 U1339 ( .A0(C1[33]), .A1(n959), .B0(n1124), .B1(n961), .C0(n1125), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N35) );
  AOI22XL U1340 ( .A0(PLAINTEXT[33]), .A1(n963), .B0(n964), .B1(n1126), .Y(
        n1125) );
  CLKINVX1 U1341 ( .A(n1127), .Y(n1126) );
  OAI221X1 U1342 ( .A0(n959), .A1(n1128), .B0(n1129), .B1(n961), .C0(n1130), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N34) );
  AOI22XL U1343 ( .A0(PLAINTEXT[32]), .A1(n963), .B0(n964), .B1(n1131), .Y(
        n1130) );
  CLKINVX1 U1344 ( .A(n1132), .Y(n1131) );
  CLKINVX1 U1345 ( .A(C1[32]), .Y(n1128) );
  OAI221X1 U1346 ( .A0(n959), .A1(n1133), .B0(n1134), .B1(n961), .C0(n1135), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N33) );
  AOI22XL U1347 ( .A0(PLAINTEXT[31]), .A1(n963), .B0(n964), .B1(n1136), .Y(
        n1135) );
  CLKINVX1 U1348 ( .A(n1137), .Y(n1136) );
  OAI221X1 U1349 ( .A0(C1[30]), .A1(n959), .B0(n1138), .B1(n961), .C0(n1139), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N32) );
  AOI22XL U1350 ( .A0(PLAINTEXT[30]), .A1(n963), .B0(n1140), .B1(n964), .Y(
        n1139) );
  OAI221X1 U1351 ( .A0(n959), .A1(n1141), .B0(n1142), .B1(n961), .C0(n1143), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N31) );
  AOI22XL U1352 ( .A0(PLAINTEXT[29]), .A1(n963), .B0(n964), .B1(n1144), .Y(
        n1143) );
  CLKINVX1 U1353 ( .A(n1145), .Y(n1144) );
  OAI221X1 U1354 ( .A0(C1[28]), .A1(n959), .B0(n1146), .B1(n961), .C0(n1147), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N30) );
  AOI22XL U1355 ( .A0(PLAINTEXT[28]), .A1(n963), .B0(n964), .B1(n1148), .Y(
        n1147) );
  CLKINVX1 U1356 ( .A(n1149), .Y(n1148) );
  OAI221X1 U1357 ( .A0(n959), .A1(n1150), .B0(n1151), .B1(n961), .C0(n1152), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N3) );
  AOI22XL U1358 ( .A0(PLAINTEXT[1]), .A1(n963), .B0(n964), .B1(n1153), .Y(
        n1152) );
  OAI221X1 U1359 ( .A0(C1[27]), .A1(n959), .B0(n1154), .B1(n961), .C0(n1155), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N29) );
  AOI22XL U1360 ( .A0(PLAINTEXT[27]), .A1(n963), .B0(n964), .B1(n1156), .Y(
        n1155) );
  CLKINVX1 U1361 ( .A(n1157), .Y(n1156) );
  OAI221X1 U1362 ( .A0(n959), .A1(n1158), .B0(n961), .B1(n1159), .C0(n1160), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N28) );
  AOI22XL U1363 ( .A0(PLAINTEXT[26]), .A1(n963), .B0(n964), .B1(n1161), .Y(
        n1160) );
  CLKINVX1 U1364 ( .A(n1162), .Y(n1161) );
  CLKINVX1 U1365 ( .A(C1[26]), .Y(n1158) );
  OAI221X1 U1366 ( .A0(C1[25]), .A1(n959), .B0(n1163), .B1(n961), .C0(n1164), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N27) );
  AOI22XL U1367 ( .A0(PLAINTEXT[25]), .A1(n963), .B0(n964), .B1(n1165), .Y(
        n1164) );
  CLKINVX1 U1368 ( .A(n1166), .Y(n1165) );
  OAI221X1 U1369 ( .A0(C1[24]), .A1(n959), .B0(n961), .B1(n1167), .C0(n1168), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N26) );
  AOI22XL U1370 ( .A0(PLAINTEXT[24]), .A1(n963), .B0(n964), .B1(n1169), .Y(
        n1168) );
  CLKINVX1 U1371 ( .A(n1170), .Y(n1169) );
  OAI221X1 U1372 ( .A0(n959), .A1(n1171), .B0(n1172), .B1(n961), .C0(n1173), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N25) );
  AOI22XL U1373 ( .A0(PLAINTEXT[23]), .A1(n963), .B0(n964), .B1(n1174), .Y(
        n1173) );
  CLKINVX1 U1374 ( .A(n1175), .Y(n1174) );
  OAI221X1 U1375 ( .A0(C1[22]), .A1(n959), .B0(n1176), .B1(n961), .C0(n1177), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N24) );
  AOI22XL U1376 ( .A0(PLAINTEXT[22]), .A1(n963), .B0(n964), .B1(n1178), .Y(
        n1177) );
  CLKINVX1 U1377 ( .A(n1179), .Y(n1178) );
  OAI221X1 U1378 ( .A0(C1[21]), .A1(n959), .B0(n961), .B1(n1180), .C0(n1181), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N23) );
  AOI22XL U1379 ( .A0(PLAINTEXT[21]), .A1(n963), .B0(n964), .B1(n1182), .Y(
        n1181) );
  CLKINVX1 U1380 ( .A(n1183), .Y(n1182) );
  OAI221X1 U1381 ( .A0(C1[20]), .A1(n959), .B0(n1184), .B1(n961), .C0(n1185), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N22) );
  AOI22XL U1382 ( .A0(PLAINTEXT[20]), .A1(n963), .B0(n964), .B1(n1186), .Y(
        n1185) );
  CLKINVX1 U1383 ( .A(n1187), .Y(n1186) );
  OAI221X1 U1384 ( .A0(C1[19]), .A1(n959), .B0(n1188), .B1(n961), .C0(n1189), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N21) );
  AOI22XL U1385 ( .A0(PLAINTEXT[19]), .A1(n963), .B0(n964), .B1(n1190), .Y(
        n1189) );
  CLKINVX1 U1386 ( .A(n1191), .Y(n1190) );
  OAI221X1 U1387 ( .A0(C1[18]), .A1(n959), .B0(n1192), .B1(n961), .C0(n1193), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N20) );
  AOI22XL U1388 ( .A0(PLAINTEXT[18]), .A1(n963), .B0(n964), .B1(n1194), .Y(
        n1193) );
  CLKINVX1 U1389 ( .A(n1195), .Y(n1194) );
  OAI221X1 U1390 ( .A0(C1[0]), .A1(n959), .B0(n1196), .B1(n961), .C0(n1197), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N2) );
  AOI22XL U1391 ( .A0(PLAINTEXT[0]), .A1(n963), .B0(n964), .B1(n1198), .Y(
        n1197) );
  CLKINVX1 U1392 ( .A(n1199), .Y(n1198) );
  OAI221X1 U1393 ( .A0(C1[17]), .A1(n959), .B0(n1200), .B1(n961), .C0(n1201), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N19) );
  AOI22XL U1394 ( .A0(PLAINTEXT[17]), .A1(n963), .B0(n964), .B1(n1202), .Y(
        n1201) );
  CLKINVX1 U1395 ( .A(n1203), .Y(n1202) );
  OAI221X1 U1396 ( .A0(C1[16]), .A1(n959), .B0(n1204), .B1(n961), .C0(n1205), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N18) );
  AOI22XL U1397 ( .A0(PLAINTEXT[16]), .A1(n963), .B0(n964), .B1(n1206), .Y(
        n1205) );
  CLKINVX1 U1398 ( .A(n1207), .Y(n1206) );
  OAI221X1 U1399 ( .A0(C1[15]), .A1(n959), .B0(n961), .B1(n1208), .C0(n1209), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N17) );
  AOI22XL U1400 ( .A0(PLAINTEXT[15]), .A1(n963), .B0(n964), .B1(n1210), .Y(
        n1209) );
  CLKINVX1 U1401 ( .A(n1211), .Y(n1210) );
  CLKINVX1 U1402 ( .A(n1212), .Y(n1208) );
  OAI221X1 U1403 ( .A0(C1[14]), .A1(n959), .B0(n1213), .B1(n961), .C0(n1214), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N16) );
  AOI22XL U1404 ( .A0(PLAINTEXT[14]), .A1(n963), .B0(n964), .B1(n1215), .Y(
        n1214) );
  CLKINVX1 U1405 ( .A(n1216), .Y(n1215) );
  OAI221X1 U1406 ( .A0(C1[13]), .A1(n959), .B0(n1217), .B1(n961), .C0(n1218), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N15) );
  AOI22XL U1407 ( .A0(PLAINTEXT[13]), .A1(n963), .B0(n964), .B1(n1219), .Y(
        n1218) );
  OAI221X1 U1408 ( .A0(n959), .A1(n1220), .B0(n1221), .B1(n961), .C0(n1222), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N14) );
  AOI22XL U1409 ( .A0(PLAINTEXT[12]), .A1(n963), .B0(n964), .B1(n1223), .Y(
        n1222) );
  CLKINVX1 U1410 ( .A(n1224), .Y(n1223) );
  OAI221X1 U1411 ( .A0(C1[11]), .A1(n959), .B0(n1225), .B1(n961), .C0(n1226), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N13) );
  AOI22XL U1412 ( .A0(PLAINTEXT[11]), .A1(n963), .B0(n964), .B1(n1227), .Y(
        n1226) );
  CLKINVX1 U1413 ( .A(n1228), .Y(n1227) );
  OAI221X1 U1414 ( .A0(C1[10]), .A1(n959), .B0(n1229), .B1(n961), .C0(n1230), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N12) );
  AOI22XL U1415 ( .A0(PLAINTEXT[10]), .A1(n963), .B0(n964), .B1(n1231), .Y(
        n1230) );
  CLKINVX1 U1416 ( .A(n1232), .Y(n1231) );
  OAI221X1 U1417 ( .A0(n959), .A1(n1233), .B0(n1234), .B1(n961), .C0(n1235), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N11) );
  AOI22XL U1418 ( .A0(PLAINTEXT[9]), .A1(n963), .B0(n964), .B1(n1236), .Y(
        n1235) );
  OAI221X1 U1419 ( .A0(n959), .A1(n1237), .B0(n1238), .B1(n961), .C0(n1239), 
        .Y(Inst_forkAE_REG_INTERNAL_STATE_N10) );
  AOI22XL U1420 ( .A0(PLAINTEXT[8]), .A1(n963), .B0(n964), .B1(n1240), .Y(
        n1239) );
  CLKINVX1 U1421 ( .A(n1241), .Y(n1240) );
  CLKINVX1 U1422 ( .A(C1[8]), .Y(n1237) );
  CLKNAND2X2 U1423 ( .A(n1242), .B(n1244), .Y(n959) );
  CLKNAND2X2 U1424 ( .A(n1244), .B(n949), .Y(n1242) );
  OAI221X1 U1425 ( .A0(n966), .A1(n1245), .B0(n1246), .B1(n1247), .C0(n1248), 
        .Y(Inst_forkAE_L_N9) );
  AOI22XL U1426 ( .A0(n1249), .A1(n1250), .B0(C1[7]), .B1(n135), .Y(n1248) );
  OAI221X1 U1427 ( .A0(n971), .A1(n1245), .B0(n968), .B1(n1247), .C0(n1252), 
        .Y(Inst_forkAE_L_N8) );
  AOI22XL U1428 ( .A0(n1249), .A1(n1253), .B0(n135), .B1(C1[6]), .Y(n1252) );
  OAI221X1 U1429 ( .A0(n1254), .A1(n1245), .B0(n973), .B1(n1247), .C0(n1255), 
        .Y(Inst_forkAE_L_N7) );
  AOI22XL U1430 ( .A0(n1249), .A1(n1256), .B0(n135), .B1(C1[5]), .Y(n1255) );
  OAI221X1 U1431 ( .A0(n1257), .A1(n1258), .B0(n1259), .B1(n1245), .C0(n1260), 
        .Y(Inst_forkAE_L_N65) );
  AOI2BB2X1 U1432 ( .B0(n135), .B1(C1[63]), .A0N(n1247), .A1N(n977), .Y(n1260)
         );
  XOR2X1 U1433 ( .A(n1212), .B(n1261), .Y(n977) );
  XNOR2X1 U1434 ( .A(n1262), .B(n1263), .Y(n1258) );
  OAI221X1 U1435 ( .A0(n1264), .A1(n1257), .B0(n984), .B1(n1245), .C0(n1265), 
        .Y(Inst_forkAE_L_N64) );
  AOI2BB2X1 U1436 ( .B0(n135), .B1(C1[62]), .A0N(n1247), .A1N(n981), .Y(n1265)
         );
  XNOR2X1 U1437 ( .A(n1213), .B(n1266), .Y(n981) );
  XNOR2X1 U1438 ( .A(n1267), .B(n1268), .Y(n1264) );
  OAI221X1 U1439 ( .A0(n1269), .A1(n1257), .B0(n989), .B1(n1245), .C0(n1270), 
        .Y(Inst_forkAE_L_N63) );
  AOI2BB2X1 U1440 ( .B0(n135), .B1(C1[61]), .A0N(n1247), .A1N(n986), .Y(n1270)
         );
  XOR2X1 U1441 ( .A(n1217), .B(n1271), .Y(n986) );
  XOR2X1 U1442 ( .A(n1272), .B(n1273), .Y(n1271) );
  NAND2BX1 U1443 ( .AN(C0[9]), .B(n1261), .Y(n1273) );
  CLKINVX1 U1444 ( .A(C0[10]), .Y(n1272) );
  CLKINVX1 U1445 ( .A(n1274), .Y(n1217) );
  XNOR2X1 U1446 ( .A(n1275), .B(n1276), .Y(n1269) );
  XNOR2X1 U1447 ( .A(C1[10]), .B(n1277), .Y(n1276) );
  CLKNAND2X2 U1448 ( .A(n1262), .B(n1233), .Y(n1277) );
  CLKINVX1 U1449 ( .A(C1[9]), .Y(n1233) );
  OAI221X1 U1450 ( .A0(n1257), .A1(n1278), .B0(n1279), .B1(n1245), .C0(n1280), 
        .Y(Inst_forkAE_L_N62) );
  AOI22XL U1451 ( .A0(n990), .A1(n1281), .B0(C1[60]), .B1(n135), .Y(n1280) );
  XOR2X1 U1452 ( .A(n1221), .B(n1282), .Y(n990) );
  XNOR2X1 U1453 ( .A(C0[9]), .B(n1283), .Y(n1282) );
  CLKNAND2X2 U1454 ( .A(n1266), .B(n1261), .Y(n1283) );
  XNOR2X1 U1455 ( .A(C0[8]), .B(n1284), .Y(n1261) );
  NOR2X1 U1456 ( .A(C0[10]), .B(C0[11]), .Y(n1284) );
  XNOR2X1 U1457 ( .A(C0[11]), .B(n1285), .Y(n1266) );
  NOR2X1 U1458 ( .A(C0[10]), .B(C0[9]), .Y(n1285) );
  CLKINVX1 U1459 ( .A(n992), .Y(n1279) );
  XOR2X1 U1460 ( .A(n1286), .B(n1287), .Y(n992) );
  CLKNAND2X2 U1461 ( .A(n984), .B(n1259), .Y(n1286) );
  CLKINVX1 U1462 ( .A(n979), .Y(n1259) );
  XOR2X1 U1463 ( .A(n1288), .B(n1289), .Y(n979) );
  CLKNAND2X2 U1464 ( .A(n984), .B(n989), .Y(n1288) );
  XOR2X1 U1465 ( .A(n1290), .B(n1291), .Y(n984) );
  XOR2X1 U1466 ( .A(C0[45]), .B(n1292), .Y(n1291) );
  XOR2X1 U1467 ( .A(Inst_forkAE_KEY_INVERSE[153]), .B(Inst_forkAE_CONST_ENC_2_), .Y(n1292) );
  XOR2X1 U1468 ( .A(n1293), .B(n1294), .Y(n1290) );
  CLKNAND2X2 U1469 ( .A(n989), .B(n1287), .Y(n1293) );
  XOR2X1 U1470 ( .A(n1295), .B(n1296), .Y(n989) );
  XOR2X1 U1471 ( .A(C0[44]), .B(n1297), .Y(n1296) );
  XOR2X1 U1472 ( .A(Inst_forkAE_KEY_INVERSE[152]), .B(Inst_forkAE_CONST_ENC_1_), .Y(n1297) );
  XOR2X1 U1473 ( .A(n1298), .B(n1299), .Y(n1295) );
  CLKNAND2X2 U1474 ( .A(n1289), .B(n1287), .Y(n1298) );
  XNOR2X1 U1475 ( .A(n1300), .B(n1301), .Y(n1287) );
  XOR2X1 U1476 ( .A(n180), .B(Inst_forkAE_KEY_INVERSE[155]), .Y(n1301) );
  XOR2X1 U1477 ( .A(n1302), .B(n1303), .Y(n1300) );
  XNOR2X1 U1478 ( .A(n1304), .B(n1305), .Y(n1289) );
  XOR2X1 U1479 ( .A(n179), .B(Inst_forkAE_KEY_INVERSE[154]), .Y(n1305) );
  XNOR2X1 U1480 ( .A(C0[46]), .B(n1306), .Y(n1304) );
  XOR2X1 U1481 ( .A(n1307), .B(n1308), .Y(n1278) );
  XOR2X1 U1482 ( .A(n1309), .B(C1[9]), .Y(n1308) );
  NAND2BX1 U1483 ( .AN(n1268), .B(n1262), .Y(n1309) );
  XNOR2X1 U1484 ( .A(C1[8]), .B(n1310), .Y(n1262) );
  NOR2X1 U1485 ( .A(C1[10]), .B(C1[11]), .Y(n1310) );
  XOR2X1 U1486 ( .A(C1[11]), .B(n1311), .Y(n1268) );
  NOR2X1 U1487 ( .A(C1[10]), .B(C1[9]), .Y(n1311) );
  OAI221X1 U1488 ( .A0(n1312), .A1(n1257), .B0(n997), .B1(n1245), .C0(n1313), 
        .Y(Inst_forkAE_L_N61) );
  AOI2BB2X1 U1489 ( .B0(n135), .B1(C1[59]), .A0N(n1247), .A1N(n994), .Y(n1313)
         );
  XNOR2X1 U1490 ( .A(n1225), .B(n1314), .Y(n994) );
  XOR2X1 U1491 ( .A(n1315), .B(n1316), .Y(n1312) );
  OAI221X1 U1492 ( .A0(n1317), .A1(n1257), .B0(n1002), .B1(n1245), .C0(n1318), 
        .Y(Inst_forkAE_L_N60) );
  AOI2BB2X1 U1493 ( .B0(n135), .B1(C1[58]), .A0N(n1247), .A1N(n999), .Y(n1318)
         );
  XNOR2X1 U1494 ( .A(n1229), .B(n1319), .Y(n999) );
  CLKINVX1 U1495 ( .A(n1320), .Y(n1229) );
  XNOR2X1 U1496 ( .A(n1321), .B(n1322), .Y(n1317) );
  OAI221X1 U1497 ( .A0(n1007), .A1(n1245), .B0(n1004), .B1(n1247), .C0(n1323), 
        .Y(Inst_forkAE_L_N6) );
  AOI22XL U1498 ( .A0(n1249), .A1(n1324), .B0(n135), .B1(C1[4]), .Y(n1323) );
  XOR2X1 U1499 ( .A(n1325), .B(n1326), .Y(n1007) );
  CLKNAND2X2 U1500 ( .A(n966), .B(n971), .Y(n1325) );
  XOR2X1 U1501 ( .A(n1327), .B(n1328), .Y(n966) );
  CLKNAND2X2 U1502 ( .A(n971), .B(n1254), .Y(n1327) );
  XOR2X1 U1503 ( .A(n1329), .B(n1330), .Y(n971) );
  XOR2X1 U1504 ( .A(C0[9]), .B(C0[57]), .Y(n1330) );
  OR2X1 U1505 ( .A(n1326), .B(n975), .Y(n1329) );
  CLKINVX1 U1506 ( .A(n1254), .Y(n975) );
  XOR2X1 U1507 ( .A(n1331), .B(n1332), .Y(n1254) );
  NOR2X1 U1508 ( .A(n1326), .B(n1328), .Y(n1332) );
  XOR2X1 U1509 ( .A(C0[10]), .B(C0[58]), .Y(n1328) );
  XNOR2X1 U1510 ( .A(C0[56]), .B(C0[8]), .Y(n1331) );
  XOR2X1 U1511 ( .A(C0[59]), .B(C0[11]), .Y(n1326) );
  OAI221X1 U1512 ( .A0(n1333), .A1(n1257), .B0(n1011), .B1(n1245), .C0(n1334), 
        .Y(Inst_forkAE_L_N59) );
  AOI22XL U1513 ( .A0(n1008), .A1(n1281), .B0(C1[57]), .B1(n135), .Y(n1334) );
  XOR2X1 U1514 ( .A(n1234), .B(n1335), .Y(n1008) );
  XNOR2X1 U1515 ( .A(C0[6]), .B(n1336), .Y(n1335) );
  CLKNAND2X2 U1516 ( .A(n1314), .B(n1337), .Y(n1336) );
  XNOR2X1 U1517 ( .A(n1338), .B(n1339), .Y(n1333) );
  XOR2X1 U1518 ( .A(n967), .B(n1340), .Y(n1339) );
  CLKNAND2X2 U1519 ( .A(n1316), .B(n972), .Y(n1340) );
  CLKINVX1 U1520 ( .A(C1[6]), .Y(n967) );
  OAI221X1 U1521 ( .A0(n1341), .A1(n1257), .B0(n1016), .B1(n1245), .C0(n1342), 
        .Y(Inst_forkAE_L_N58) );
  AOI2BB2X1 U1522 ( .B0(n135), .B1(C1[56]), .A0N(n1247), .A1N(n1013), .Y(n1342) );
  XOR2X1 U1523 ( .A(n1238), .B(n1343), .Y(n1013) );
  XOR2X1 U1524 ( .A(n1337), .B(n1344), .Y(n1343) );
  CLKNAND2X2 U1525 ( .A(n1319), .B(n1314), .Y(n1344) );
  XNOR2X1 U1526 ( .A(C0[4]), .B(n1345), .Y(n1314) );
  NOR2X1 U1527 ( .A(C0[6]), .B(C0[7]), .Y(n1345) );
  XNOR2X1 U1528 ( .A(C0[7]), .B(n1346), .Y(n1319) );
  NOR2X1 U1529 ( .A(C0[5]), .B(C0[6]), .Y(n1346) );
  CLKINVX1 U1530 ( .A(C0[5]), .Y(n1337) );
  XNOR2X1 U1531 ( .A(n1347), .B(n1348), .Y(n1016) );
  CLKNAND2X2 U1532 ( .A(n997), .B(n1002), .Y(n1347) );
  XOR2X1 U1533 ( .A(n1349), .B(n1350), .Y(n997) );
  CLKNAND2X2 U1534 ( .A(n1002), .B(n1011), .Y(n1349) );
  XOR2X1 U1535 ( .A(n1351), .B(n1352), .Y(n1002) );
  XOR2X1 U1536 ( .A(Inst_forkAE_KEY_INVERSE[129]), .B(C0[41]), .Y(n1352) );
  XOR2X1 U1537 ( .A(n1353), .B(n1354), .Y(n1351) );
  CLKNAND2X2 U1538 ( .A(n1011), .B(n1348), .Y(n1353) );
  XOR2X1 U1539 ( .A(n1355), .B(n1356), .Y(n1011) );
  XOR2X1 U1540 ( .A(Inst_forkAE_KEY_INVERSE[128]), .B(C0[40]), .Y(n1356) );
  XOR2X1 U1541 ( .A(n1357), .B(n1358), .Y(n1355) );
  NAND2BX1 U1542 ( .AN(n1350), .B(n1348), .Y(n1357) );
  XOR2X1 U1543 ( .A(n1359), .B(n1360), .Y(n1348) );
  XNOR2X1 U1544 ( .A(Inst_forkAE_KEY_INVERSE[131]), .B(C0[43]), .Y(n1359) );
  XNOR2X1 U1545 ( .A(n1361), .B(n1362), .Y(n1350) );
  XNOR2X1 U1546 ( .A(Inst_forkAE_KEY_INVERSE[130]), .B(C0[42]), .Y(n1361) );
  XNOR2X1 U1547 ( .A(n1363), .B(n1364), .Y(n1341) );
  XOR2X1 U1548 ( .A(n972), .B(n1365), .Y(n1364) );
  NAND2BX1 U1549 ( .AN(n1322), .B(n1316), .Y(n1365) );
  XOR2X1 U1550 ( .A(n1003), .B(n1366), .Y(n1316) );
  NOR2X1 U1551 ( .A(C1[7]), .B(C1[6]), .Y(n1366) );
  CLKINVX1 U1552 ( .A(C1[4]), .Y(n1003) );
  XOR2X1 U1553 ( .A(C1[7]), .B(n1367), .Y(n1322) );
  NOR2X1 U1554 ( .A(C1[5]), .B(C1[6]), .Y(n1367) );
  CLKINVX1 U1555 ( .A(C1[5]), .Y(n972) );
  OAI221X1 U1556 ( .A0(n1368), .A1(n1257), .B0(n1021), .B1(n1245), .C0(n1369), 
        .Y(Inst_forkAE_L_N57) );
  AOI2BB2X1 U1557 ( .B0(n135), .B1(C1[55]), .A0N(n1247), .A1N(n1018), .Y(n1369) );
  XNOR2X1 U1558 ( .A(n960), .B(n1370), .Y(n1018) );
  CLKINVX1 U1559 ( .A(n1246), .Y(n960) );
  XOR2X1 U1560 ( .A(n1093), .B(n1371), .Y(n1246) );
  XOR2X1 U1561 ( .A(n1250), .B(n1372), .Y(n1368) );
  XNOR2X1 U1562 ( .A(n1373), .B(n1374), .Y(n1250) );
  OAI221X1 U1563 ( .A0(n1375), .A1(n1257), .B0(n1376), .B1(n1245), .C0(n1377), 
        .Y(Inst_forkAE_L_N56) );
  AOI22XL U1564 ( .A0(n1022), .A1(n1281), .B0(C1[54]), .B1(n135), .Y(n1377) );
  XNOR2X1 U1565 ( .A(n968), .B(n1378), .Y(n1022) );
  XOR2X1 U1566 ( .A(n1097), .B(n1379), .Y(n968) );
  CLKINVX1 U1567 ( .A(n1380), .Y(n1379) );
  XNOR2X1 U1568 ( .A(n1253), .B(n1381), .Y(n1375) );
  XOR2X1 U1569 ( .A(n1382), .B(n1383), .Y(n1253) );
  CLKINVX1 U1570 ( .A(n1384), .Y(n1383) );
  OAI221X1 U1571 ( .A0(n1385), .A1(n1257), .B0(n1029), .B1(n1245), .C0(n1386), 
        .Y(Inst_forkAE_L_N55) );
  AOI2BB2X1 U1572 ( .B0(n135), .B1(C1[53]), .A0N(n1247), .A1N(n1026), .Y(n1386) );
  XOR2X1 U1573 ( .A(n973), .B(n1387), .Y(n1026) );
  XNOR2X1 U1574 ( .A(C0[2]), .B(n1388), .Y(n1387) );
  CLKNAND2X2 U1575 ( .A(n1370), .B(n1389), .Y(n1388) );
  XNOR2X1 U1576 ( .A(n1107), .B(n1390), .Y(n973) );
  XNOR2X1 U1577 ( .A(n1256), .B(n1391), .Y(n1385) );
  XOR2X1 U1578 ( .A(n1101), .B(n1392), .Y(n1391) );
  CLKNAND2X2 U1579 ( .A(n1372), .B(n1150), .Y(n1392) );
  CLKINVX1 U1580 ( .A(C1[2]), .Y(n1101) );
  XNOR2X1 U1581 ( .A(n1393), .B(n1394), .Y(n1256) );
  CLKINVX1 U1582 ( .A(n1395), .Y(n1394) );
  OAI221X1 U1583 ( .A0(n1396), .A1(n1257), .B0(n1034), .B1(n1245), .C0(n1397), 
        .Y(Inst_forkAE_L_N54) );
  AOI2BB2X1 U1584 ( .B0(n135), .B1(C1[52]), .A0N(n1247), .A1N(n1031), .Y(n1397) );
  XOR2X1 U1585 ( .A(n1004), .B(n1398), .Y(n1031) );
  XOR2X1 U1586 ( .A(n1389), .B(n1399), .Y(n1398) );
  CLKNAND2X2 U1587 ( .A(n1378), .B(n1370), .Y(n1399) );
  XNOR2X1 U1588 ( .A(C0[0]), .B(n1400), .Y(n1370) );
  NOR2X1 U1589 ( .A(C0[2]), .B(C0[3]), .Y(n1400) );
  XNOR2X1 U1590 ( .A(C0[3]), .B(n1401), .Y(n1378) );
  NOR2X1 U1591 ( .A(C0[1]), .B(C0[2]), .Y(n1401) );
  CLKINVX1 U1592 ( .A(C0[1]), .Y(n1389) );
  XOR2X1 U1593 ( .A(n1111), .B(n1402), .Y(n1004) );
  XNOR2X1 U1594 ( .A(n1403), .B(n1404), .Y(n1034) );
  CLKNAND2X2 U1595 ( .A(n1021), .B(n1376), .Y(n1403) );
  XOR2X1 U1596 ( .A(n1405), .B(n1406), .Y(n1021) );
  CLKNAND2X2 U1597 ( .A(n1029), .B(n1376), .Y(n1405) );
  CLKINVX1 U1598 ( .A(n1024), .Y(n1376) );
  XOR2X1 U1599 ( .A(n1407), .B(n1408), .Y(n1024) );
  XOR2X1 U1600 ( .A(n1409), .B(C0[37]), .Y(n1407) );
  CLKNAND2X2 U1601 ( .A(n1029), .B(n1404), .Y(n1409) );
  XOR2X1 U1602 ( .A(n1410), .B(n1411), .Y(n1029) );
  XOR2X1 U1603 ( .A(Inst_forkAE_KEY_INVERSE[156]), .B(C0[36]), .Y(n1411) );
  XOR2X1 U1604 ( .A(n1412), .B(n1413), .Y(n1410) );
  NAND2BX1 U1605 ( .AN(n1406), .B(n1404), .Y(n1412) );
  XOR2X1 U1606 ( .A(n1414), .B(n1415), .Y(n1404) );
  XNOR2X1 U1607 ( .A(Inst_forkAE_KEY_INVERSE[159]), .B(C0[39]), .Y(n1414) );
  XNOR2X1 U1608 ( .A(n1416), .B(n1417), .Y(n1406) );
  XOR2X1 U1609 ( .A(Inst_forkAE_KEY_INVERSE[158]), .B(n1418), .Y(n1416) );
  XNOR2X1 U1610 ( .A(n1324), .B(n1419), .Y(n1396) );
  XOR2X1 U1611 ( .A(n1150), .B(n1420), .Y(n1419) );
  NAND2BX1 U1612 ( .AN(n1381), .B(n1372), .Y(n1420) );
  XNOR2X1 U1613 ( .A(C1[0]), .B(n1421), .Y(n1372) );
  NOR2X1 U1614 ( .A(C1[2]), .B(C1[3]), .Y(n1421) );
  XNOR2X1 U1615 ( .A(n1053), .B(n1422), .Y(n1381) );
  NOR2X1 U1616 ( .A(C1[1]), .B(C1[2]), .Y(n1422) );
  CLKINVX1 U1617 ( .A(C1[3]), .Y(n1053) );
  CLKINVX1 U1618 ( .A(C1[1]), .Y(n1150) );
  XOR2X1 U1619 ( .A(n1423), .B(n1424), .Y(n1324) );
  CLKINVX1 U1620 ( .A(n1425), .Y(n1424) );
  OAI221X1 U1621 ( .A0(n1426), .A1(n1257), .B0(n1038), .B1(n1245), .C0(n1427), 
        .Y(Inst_forkAE_L_N53) );
  AOI22XL U1622 ( .A0(n1035), .A1(n1281), .B0(C1[51]), .B1(n135), .Y(n1427) );
  XNOR2X1 U1623 ( .A(n1054), .B(n1428), .Y(n1035) );
  XOR2X1 U1624 ( .A(n1429), .B(n1430), .Y(n1426) );
  OAI221X1 U1625 ( .A0(n1431), .A1(n1257), .B0(n1043), .B1(n1245), .C0(n1432), 
        .Y(Inst_forkAE_L_N52) );
  AOI2BB2X1 U1626 ( .B0(n135), .B1(C1[50]), .A0N(n1247), .A1N(n1040), .Y(n1432) );
  XNOR2X1 U1627 ( .A(n1102), .B(n1433), .Y(n1040) );
  XNOR2X1 U1628 ( .A(n1434), .B(n1435), .Y(n1431) );
  OAI221X1 U1629 ( .A0(n1436), .A1(n1257), .B0(n1048), .B1(n1245), .C0(n1437), 
        .Y(Inst_forkAE_L_N51) );
  AOI2BB2X1 U1630 ( .B0(n135), .B1(C1[49]), .A0N(n1247), .A1N(n1045), .Y(n1437) );
  XOR2X1 U1631 ( .A(n1151), .B(n1438), .Y(n1045) );
  XNOR2X1 U1632 ( .A(C0[14]), .B(n1439), .Y(n1438) );
  CLKNAND2X2 U1633 ( .A(n1428), .B(n1440), .Y(n1439) );
  XNOR2X1 U1634 ( .A(n1441), .B(n1442), .Y(n1436) );
  XNOR2X1 U1635 ( .A(C1[14]), .B(n1443), .Y(n1442) );
  NAND2BX1 U1636 ( .AN(C1[13]), .B(n1430), .Y(n1443) );
  OAI221X1 U1637 ( .A0(n1444), .A1(n1257), .B0(n1052), .B1(n1245), .C0(n1445), 
        .Y(Inst_forkAE_L_N50) );
  AOI22XL U1638 ( .A0(n1049), .A1(n1281), .B0(C1[48]), .B1(n135), .Y(n1445) );
  XOR2X1 U1639 ( .A(n1196), .B(n1446), .Y(n1049) );
  XOR2X1 U1640 ( .A(n1440), .B(n1447), .Y(n1446) );
  CLKNAND2X2 U1641 ( .A(n1433), .B(n1428), .Y(n1447) );
  XNOR2X1 U1642 ( .A(C0[12]), .B(n1448), .Y(n1428) );
  NOR2X1 U1643 ( .A(C0[14]), .B(C0[15]), .Y(n1448) );
  XNOR2X1 U1644 ( .A(C0[15]), .B(n1449), .Y(n1433) );
  NOR2X1 U1645 ( .A(C0[13]), .B(C0[14]), .Y(n1449) );
  CLKINVX1 U1646 ( .A(C0[13]), .Y(n1440) );
  XNOR2X1 U1647 ( .A(n1450), .B(n1451), .Y(n1052) );
  CLKNAND2X2 U1648 ( .A(n1038), .B(n1043), .Y(n1450) );
  XOR2X1 U1649 ( .A(n1452), .B(n1453), .Y(n1038) );
  CLKNAND2X2 U1650 ( .A(n1043), .B(n1048), .Y(n1452) );
  XOR2X1 U1651 ( .A(n1454), .B(n1455), .Y(n1043) );
  XOR2X1 U1652 ( .A(Inst_forkAE_KEY_INVERSE[137]), .B(C0[33]), .Y(n1455) );
  XOR2X1 U1653 ( .A(n1456), .B(n1457), .Y(n1454) );
  CLKNAND2X2 U1654 ( .A(n1048), .B(n1451), .Y(n1456) );
  XOR2X1 U1655 ( .A(n1458), .B(n1459), .Y(n1048) );
  XOR2X1 U1656 ( .A(Inst_forkAE_KEY_INVERSE[136]), .B(C0[32]), .Y(n1459) );
  XOR2X1 U1657 ( .A(n1460), .B(n1461), .Y(n1458) );
  NAND2BX1 U1658 ( .AN(n1453), .B(n1451), .Y(n1460) );
  XOR2X1 U1659 ( .A(n1462), .B(n1463), .Y(n1451) );
  XNOR2X1 U1660 ( .A(Inst_forkAE_KEY_INVERSE[139]), .B(C0[35]), .Y(n1462) );
  XNOR2X1 U1661 ( .A(n1464), .B(n1465), .Y(n1453) );
  XNOR2X1 U1662 ( .A(Inst_forkAE_KEY_INVERSE[138]), .B(C0[34]), .Y(n1464) );
  XNOR2X1 U1663 ( .A(n1466), .B(n1467), .Y(n1444) );
  XNOR2X1 U1664 ( .A(C1[13]), .B(n1468), .Y(n1467) );
  NAND2BX1 U1665 ( .AN(n1435), .B(n1430), .Y(n1468) );
  XOR2X1 U1666 ( .A(n1220), .B(n1469), .Y(n1430) );
  NOR2X1 U1667 ( .A(C1[14]), .B(C1[15]), .Y(n1469) );
  CLKINVX1 U1668 ( .A(C1[12]), .Y(n1220) );
  XOR2X1 U1669 ( .A(C1[15]), .B(n1470), .Y(n1435) );
  NOR2X1 U1670 ( .A(C1[13]), .B(C1[14]), .Y(n1470) );
  OAI221X1 U1671 ( .A0(n1057), .A1(n1245), .B0(n1054), .B1(n1247), .C0(n1471), 
        .Y(Inst_forkAE_L_N5) );
  AOI22XL U1672 ( .A0(n1249), .A1(n1429), .B0(n135), .B1(C1[3]), .Y(n1471) );
  XNOR2X1 U1673 ( .A(n1472), .B(n1473), .Y(n1429) );
  XOR2X1 U1674 ( .A(n1474), .B(n1475), .Y(n1054) );
  OAI221X1 U1675 ( .A0(n1062), .A1(n1245), .B0(n1059), .B1(n1247), .C0(n1476), 
        .Y(Inst_forkAE_L_N49) );
  AOI22XL U1676 ( .A0(n1477), .A1(n1249), .B0(n135), .B1(C1[47]), .Y(n1476) );
  OAI221X1 U1677 ( .A0(n1478), .A1(n1245), .B0(n1064), .B1(n1247), .C0(n1479), 
        .Y(Inst_forkAE_L_N48) );
  AOI22XL U1678 ( .A0(n1249), .A1(n1480), .B0(n135), .B1(C1[46]), .Y(n1479) );
  OAI221X1 U1679 ( .A0(n1070), .A1(n1245), .B0(n1481), .B1(n1247), .C0(n1482), 
        .Y(Inst_forkAE_L_N47) );
  AOI22XL U1680 ( .A0(n1249), .A1(n1483), .B0(C1[45]), .B1(n135), .Y(n1482) );
  CLKINVX1 U1681 ( .A(n1067), .Y(n1481) );
  OAI221X1 U1682 ( .A0(n1074), .A1(n1245), .B0(n1484), .B1(n1247), .C0(n1485), 
        .Y(Inst_forkAE_L_N46) );
  AOI22XL U1683 ( .A0(n1486), .A1(n1249), .B0(C1[44]), .B1(n135), .Y(n1485) );
  CLKINVX1 U1684 ( .A(n1071), .Y(n1484) );
  XNOR2X1 U1685 ( .A(n1487), .B(n1488), .Y(n1074) );
  CLKNAND2X2 U1686 ( .A(n1062), .B(n1478), .Y(n1487) );
  XOR2X1 U1687 ( .A(n1489), .B(n1490), .Y(n1062) );
  CLKNAND2X2 U1688 ( .A(n1070), .B(n1478), .Y(n1489) );
  CLKINVX1 U1689 ( .A(n1066), .Y(n1478) );
  XOR2X1 U1690 ( .A(n1491), .B(n1492), .Y(n1066) );
  XOR2X1 U1691 ( .A(C0[25]), .B(n1493), .Y(n1492) );
  XOR2X1 U1692 ( .A(n181), .B(Inst_forkAE_KEY_INVERSE[149]), .Y(n1493) );
  XOR2X1 U1693 ( .A(n1494), .B(n1495), .Y(n1491) );
  XOR2X1 U1694 ( .A(n1496), .B(n1497), .Y(n1494) );
  CLKNAND2X2 U1695 ( .A(n1070), .B(n1488), .Y(n1496) );
  XOR2X1 U1696 ( .A(n1498), .B(n1499), .Y(n1070) );
  XOR2X1 U1697 ( .A(C0[24]), .B(n1500), .Y(n1499) );
  XOR2X1 U1698 ( .A(Inst_forkAE_KEY_INVERSE[148]), .B(Inst_forkAE_CONST_ENC_5_), .Y(n1500) );
  XOR2X1 U1699 ( .A(n1501), .B(n1502), .Y(n1498) );
  CLKINVX1 U1700 ( .A(n1503), .Y(n1502) );
  XOR2X1 U1701 ( .A(n1504), .B(n1505), .Y(n1501) );
  NAND2BX1 U1702 ( .AN(n1490), .B(n1488), .Y(n1504) );
  XNOR2X1 U1703 ( .A(n1506), .B(n1507), .Y(n1488) );
  XOR2X1 U1704 ( .A(n1508), .B(C0[27]), .Y(n1506) );
  XNOR2X1 U1705 ( .A(n1509), .B(n1510), .Y(n1490) );
  XOR2X1 U1706 ( .A(n1511), .B(n1512), .Y(n1510) );
  XNOR2X1 U1707 ( .A(C0[26]), .B(n1513), .Y(n1509) );
  XOR2X1 U1708 ( .A(Inst_forkAE_KEY_INVERSE[150]), .B(Inst_forkAE_CONST_DEC_6_), .Y(n1513) );
  OAI221X1 U1709 ( .A0(n1079), .A1(n1245), .B0(n1076), .B1(n1247), .C0(n1514), 
        .Y(Inst_forkAE_L_N45) );
  AOI22XL U1710 ( .A0(n1249), .A1(n1515), .B0(n135), .B1(C1[43]), .Y(n1514) );
  OAI221X1 U1711 ( .A0(n1083), .A1(n1245), .B0(n1516), .B1(n1247), .C0(n1517), 
        .Y(Inst_forkAE_L_N44) );
  AOI22XL U1712 ( .A0(n1249), .A1(n1518), .B0(C1[42]), .B1(n135), .Y(n1517) );
  CLKINVX1 U1713 ( .A(n1080), .Y(n1516) );
  OAI221X1 U1714 ( .A0(n1087), .A1(n1245), .B0(n1519), .B1(n1247), .C0(n1520), 
        .Y(Inst_forkAE_L_N43) );
  AOI22XL U1715 ( .A0(n1249), .A1(n1521), .B0(C1[41]), .B1(n135), .Y(n1520) );
  CLKINVX1 U1716 ( .A(n1084), .Y(n1519) );
  OAI221X1 U1717 ( .A0(n1092), .A1(n1245), .B0(n1089), .B1(n1247), .C0(n1522), 
        .Y(Inst_forkAE_L_N42) );
  AOI22XL U1718 ( .A0(n1249), .A1(n1523), .B0(n135), .B1(C1[40]), .Y(n1522) );
  XNOR2X1 U1719 ( .A(n1524), .B(n1525), .Y(n1092) );
  CLKNAND2X2 U1720 ( .A(n1079), .B(n1083), .Y(n1524) );
  XOR2X1 U1721 ( .A(n1526), .B(n1527), .Y(n1079) );
  CLKNAND2X2 U1722 ( .A(n1083), .B(n1087), .Y(n1526) );
  XOR2X1 U1723 ( .A(n1528), .B(n1529), .Y(n1083) );
  XOR2X1 U1724 ( .A(n1530), .B(n1531), .Y(n1529) );
  XOR2X1 U1725 ( .A(n1532), .B(n1533), .Y(n1528) );
  XOR2X1 U1726 ( .A(Inst_forkAE_KEY_INVERSE[133]), .B(C0[21]), .Y(n1533) );
  CLKNAND2X2 U1727 ( .A(n1087), .B(n1525), .Y(n1532) );
  XOR2X1 U1728 ( .A(n1534), .B(n1535), .Y(n1087) );
  XOR2X1 U1729 ( .A(n1536), .B(n1537), .Y(n1535) );
  CLKINVX1 U1730 ( .A(n1538), .Y(n1536) );
  XOR2X1 U1731 ( .A(n1539), .B(C0[20]), .Y(n1534) );
  NAND2BX1 U1732 ( .AN(n1527), .B(n1525), .Y(n1539) );
  XNOR2X1 U1733 ( .A(n1540), .B(n1541), .Y(n1525) );
  XOR2X1 U1734 ( .A(n1542), .B(C0[23]), .Y(n1540) );
  XNOR2X1 U1735 ( .A(n1543), .B(n1544), .Y(n1527) );
  XNOR2X1 U1736 ( .A(C0[22]), .B(n1545), .Y(n1543) );
  OAI221X1 U1737 ( .A0(n1096), .A1(n1245), .B0(n1546), .B1(n1247), .C0(n1547), 
        .Y(Inst_forkAE_L_N41) );
  AOI22XL U1738 ( .A0(n1249), .A1(n1373), .B0(C1[39]), .B1(n135), .Y(n1547) );
  XNOR2X1 U1739 ( .A(n1548), .B(n1549), .Y(n1373) );
  XOR2X1 U1740 ( .A(Inst_forkAE_KEY_INVERSE[114]), .B(n1550), .Y(n1549) );
  XOR2X1 U1741 ( .A(Inst_forkAE_KEY_INVERSE[48]), .B(
        Inst_forkAE_KEY_INVERSE[179]), .Y(n1550) );
  XNOR2X1 U1742 ( .A(n1551), .B(n1552), .Y(n1548) );
  CLKINVX1 U1743 ( .A(n1093), .Y(n1546) );
  XNOR2X1 U1744 ( .A(n1553), .B(n1554), .Y(n1093) );
  XNOR2X1 U1745 ( .A(Inst_forkAE_KEY_INVERSE[159]), .B(n1415), .Y(n1553) );
  XOR2X1 U1746 ( .A(Inst_forkAE_CURRENT_KEY_55_), .B(
        Inst_forkAE_KEY_INVERSE[94]), .Y(n1415) );
  OAI221X1 U1747 ( .A0(n1100), .A1(n1245), .B0(n1555), .B1(n1247), .C0(n1556), 
        .Y(Inst_forkAE_L_N40) );
  AOI22XL U1748 ( .A0(n1249), .A1(n1382), .B0(C1[38]), .B1(n135), .Y(n1556) );
  XNOR2X1 U1749 ( .A(n1557), .B(n1558), .Y(n1382) );
  XOR2X1 U1750 ( .A(Inst_forkAE_KEY_INVERSE[178]), .B(n1559), .Y(n1558) );
  XOR2X1 U1751 ( .A(Inst_forkAE_KEY_INVERSE[51]), .B(
        Inst_forkAE_KEY_INVERSE[50]), .Y(n1559) );
  XNOR2X1 U1752 ( .A(n1551), .B(n1560), .Y(n1557) );
  XOR2X1 U1753 ( .A(n696), .B(n873), .Y(n1551) );
  CLKINVX1 U1754 ( .A(Inst_forkAE_KEY_INVERSE[113]), .Y(n696) );
  CLKINVX1 U1755 ( .A(n1097), .Y(n1555) );
  XNOR2X1 U1756 ( .A(n1561), .B(n1562), .Y(n1097) );
  XNOR2X1 U1757 ( .A(Inst_forkAE_KEY_INVERSE[158]), .B(n1417), .Y(n1561) );
  XOR2X1 U1758 ( .A(Inst_forkAE_KEY_INVERSE[31]), .B(
        Inst_forkAE_KEY_INVERSE[93]), .Y(n1417) );
  OAI221X1 U1759 ( .A0(n1105), .A1(n1245), .B0(n1102), .B1(n1247), .C0(n1563), 
        .Y(Inst_forkAE_L_N4) );
  AOI22XL U1760 ( .A0(n1249), .A1(n1434), .B0(n135), .B1(C1[2]), .Y(n1563) );
  XOR2X1 U1761 ( .A(n1564), .B(n1565), .Y(n1434) );
  XOR2X1 U1762 ( .A(n1120), .B(n1566), .Y(n1102) );
  CLKINVX1 U1763 ( .A(n1567), .Y(n1566) );
  OAI221X1 U1764 ( .A0(n1110), .A1(n1245), .B0(n1107), .B1(n1247), .C0(n1568), 
        .Y(Inst_forkAE_L_N39) );
  AOI22XL U1765 ( .A0(n1393), .A1(n1249), .B0(n135), .B1(C1[37]), .Y(n1568) );
  XOR2X1 U1766 ( .A(n1569), .B(n1570), .Y(n1393) );
  XOR2X1 U1767 ( .A(n507), .B(n873), .Y(n1570) );
  XOR2X1 U1768 ( .A(Inst_forkAE_KEY_INVERSE[112]), .B(
        Inst_forkAE_KEY_INVERSE[115]), .Y(n873) );
  XOR2X1 U1769 ( .A(n530), .B(n520), .Y(n507) );
  CLKINVX1 U1770 ( .A(Inst_forkAE_KEY_INVERSE[50]), .Y(n520) );
  CLKINVX1 U1771 ( .A(Inst_forkAE_KEY_INVERSE[49]), .Y(n530) );
  XOR2X1 U1772 ( .A(n1571), .B(n1572), .Y(n1569) );
  XOR2X1 U1773 ( .A(Inst_forkAE_KEY_INVERSE[177]), .B(C1[54]), .Y(n1572) );
  CLKNAND2X2 U1774 ( .A(n1552), .B(n1025), .Y(n1571) );
  CLKINVX1 U1775 ( .A(C1[53]), .Y(n1025) );
  XNOR2X1 U1776 ( .A(n1573), .B(n1408), .Y(n1107) );
  XOR2X1 U1777 ( .A(Inst_forkAE_KEY_INVERSE[157]), .B(n1574), .Y(n1408) );
  XOR2X1 U1778 ( .A(Inst_forkAE_KEY_INVERSE[92]), .B(
        Inst_forkAE_KEY_INVERSE[30]), .Y(n1574) );
  XOR2X1 U1779 ( .A(n1575), .B(C0[54]), .Y(n1573) );
  NAND2BX1 U1780 ( .AN(C0[53]), .B(n1554), .Y(n1575) );
  OAI221X1 U1781 ( .A0(n1114), .A1(n1245), .B0(n1576), .B1(n1247), .C0(n1577), 
        .Y(Inst_forkAE_L_N38) );
  AOI22XL U1782 ( .A0(n1249), .A1(n1423), .B0(C1[36]), .B1(n135), .Y(n1577) );
  XNOR2X1 U1783 ( .A(n1578), .B(n1579), .Y(n1423) );
  XOR2X1 U1784 ( .A(Inst_forkAE_KEY_INVERSE[176]), .B(n1580), .Y(n1579) );
  XOR2X1 U1785 ( .A(Inst_forkAE_KEY_INVERSE[49]), .B(
        Inst_forkAE_KEY_INVERSE[48]), .Y(n1580) );
  XOR2X1 U1786 ( .A(n1581), .B(n1582), .Y(n1578) );
  XOR2X1 U1787 ( .A(Inst_forkAE_KEY_INVERSE[115]), .B(C1[53]), .Y(n1582) );
  CLKNAND2X2 U1788 ( .A(n1560), .B(n1552), .Y(n1581) );
  XNOR2X1 U1789 ( .A(C1[52]), .B(n1583), .Y(n1552) );
  NOR2X1 U1790 ( .A(C1[54]), .B(C1[55]), .Y(n1583) );
  XNOR2X1 U1791 ( .A(C1[55]), .B(n1584), .Y(n1560) );
  NOR2X1 U1792 ( .A(C1[54]), .B(C1[53]), .Y(n1584) );
  CLKINVX1 U1793 ( .A(n1111), .Y(n1576) );
  XOR2X1 U1794 ( .A(n1585), .B(n1586), .Y(n1111) );
  XOR2X1 U1795 ( .A(Inst_forkAE_KEY_INVERSE[156]), .B(C0[53]), .Y(n1586) );
  XOR2X1 U1796 ( .A(n1587), .B(n1413), .Y(n1585) );
  XOR2X1 U1797 ( .A(Inst_forkAE_CURRENT_KEY_116_), .B(
        Inst_forkAE_KEY_INVERSE[29]), .Y(n1413) );
  CLKNAND2X2 U1798 ( .A(n1562), .B(n1554), .Y(n1587) );
  XNOR2X1 U1799 ( .A(C0[52]), .B(n1588), .Y(n1554) );
  NOR2X1 U1800 ( .A(C0[54]), .B(C0[55]), .Y(n1588) );
  XNOR2X1 U1801 ( .A(C0[55]), .B(n1589), .Y(n1562) );
  NOR2X1 U1802 ( .A(C0[53]), .B(C0[54]), .Y(n1589) );
  XNOR2X1 U1803 ( .A(n1590), .B(n1591), .Y(n1114) );
  CLKNAND2X2 U1804 ( .A(n1096), .B(n1100), .Y(n1590) );
  XOR2X1 U1805 ( .A(n1592), .B(n1593), .Y(n1096) );
  CLKNAND2X2 U1806 ( .A(n1100), .B(n1110), .Y(n1592) );
  XOR2X1 U1807 ( .A(n1594), .B(n1595), .Y(n1100) );
  XOR2X1 U1808 ( .A(n1596), .B(n1597), .Y(n1595) );
  XOR2X1 U1809 ( .A(n1598), .B(C0[17]), .Y(n1594) );
  CLKNAND2X2 U1810 ( .A(n1110), .B(n1591), .Y(n1598) );
  XOR2X1 U1811 ( .A(n1599), .B(n1600), .Y(n1110) );
  XOR2X1 U1812 ( .A(n1601), .B(n1602), .Y(n1600) );
  XOR2X1 U1813 ( .A(n1603), .B(C0[16]), .Y(n1599) );
  NAND2BX1 U1814 ( .AN(n1593), .B(n1591), .Y(n1603) );
  XNOR2X1 U1815 ( .A(n1604), .B(n1605), .Y(n1591) );
  XOR2X1 U1816 ( .A(n1606), .B(C0[19]), .Y(n1604) );
  XNOR2X1 U1817 ( .A(n1607), .B(n1608), .Y(n1593) );
  XNOR2X1 U1818 ( .A(C0[18]), .B(n1609), .Y(n1607) );
  OAI221X1 U1819 ( .A0(n1118), .A1(n1245), .B0(n1474), .B1(n1247), .C0(n1610), 
        .Y(Inst_forkAE_L_N37) );
  AOI22XL U1820 ( .A0(n1249), .A1(n1472), .B0(C1[35]), .B1(n135), .Y(n1610) );
  XNOR2X1 U1821 ( .A(n1611), .B(n1612), .Y(n1472) );
  XOR2X1 U1822 ( .A(Inst_forkAE_KEY_INVERSE[118]), .B(n1613), .Y(n1612) );
  XOR2X1 U1823 ( .A(Inst_forkAE_KEY_INVERSE[52]), .B(
        Inst_forkAE_KEY_INVERSE[183]), .Y(n1613) );
  XNOR2X1 U1824 ( .A(n1614), .B(n1615), .Y(n1611) );
  CLKINVX1 U1825 ( .A(n1115), .Y(n1474) );
  XNOR2X1 U1826 ( .A(n1616), .B(n1617), .Y(n1115) );
  XNOR2X1 U1827 ( .A(Inst_forkAE_KEY_INVERSE[139]), .B(n1463), .Y(n1616) );
  XOR2X1 U1828 ( .A(Inst_forkAE_CURRENT_KEY_51_), .B(
        Inst_forkAE_KEY_INVERSE[74]), .Y(n1463) );
  OAI221X1 U1829 ( .A0(n1123), .A1(n1245), .B0(n1120), .B1(n1247), .C0(n1618), 
        .Y(Inst_forkAE_L_N36) );
  AOI22XL U1830 ( .A0(n1249), .A1(n1564), .B0(n135), .B1(C1[34]), .Y(n1618) );
  XNOR2X1 U1831 ( .A(n1619), .B(n1620), .Y(n1564) );
  XOR2X1 U1832 ( .A(Inst_forkAE_KEY_INVERSE[182]), .B(n1621), .Y(n1620) );
  XOR2X1 U1833 ( .A(Inst_forkAE_KEY_INVERSE[55]), .B(
        Inst_forkAE_KEY_INVERSE[54]), .Y(n1621) );
  XNOR2X1 U1834 ( .A(n1614), .B(n1622), .Y(n1619) );
  XOR2X1 U1835 ( .A(n672), .B(n899), .Y(n1614) );
  CLKINVX1 U1836 ( .A(Inst_forkAE_KEY_INVERSE[117]), .Y(n672) );
  XNOR2X1 U1837 ( .A(n1623), .B(n1624), .Y(n1120) );
  XNOR2X1 U1838 ( .A(Inst_forkAE_KEY_INVERSE[138]), .B(n1465), .Y(n1623) );
  XOR2X1 U1839 ( .A(Inst_forkAE_KEY_INVERSE[11]), .B(
        Inst_forkAE_KEY_INVERSE[73]), .Y(n1465) );
  OAI221X1 U1840 ( .A0(n1127), .A1(n1245), .B0(n1625), .B1(n1247), .C0(n1626), 
        .Y(Inst_forkAE_L_N35) );
  AOI22XL U1841 ( .A0(n1249), .A1(n1627), .B0(C1[33]), .B1(n135), .Y(n1626) );
  CLKINVX1 U1842 ( .A(n1124), .Y(n1625) );
  OAI221X1 U1843 ( .A0(n1132), .A1(n1245), .B0(n1129), .B1(n1247), .C0(n1628), 
        .Y(Inst_forkAE_L_N34) );
  AOI22XL U1844 ( .A0(n1249), .A1(n1629), .B0(n135), .B1(C1[32]), .Y(n1628) );
  XNOR2X1 U1845 ( .A(n1630), .B(n1631), .Y(n1132) );
  CLKNAND2X2 U1846 ( .A(n1118), .B(n1123), .Y(n1630) );
  XOR2X1 U1847 ( .A(n1632), .B(n1633), .Y(n1118) );
  CLKNAND2X2 U1848 ( .A(n1123), .B(n1127), .Y(n1632) );
  XOR2X1 U1849 ( .A(n1634), .B(n1635), .Y(n1123) );
  XOR2X1 U1850 ( .A(n1636), .B(n1637), .Y(n1635) );
  XOR2X1 U1851 ( .A(n1638), .B(C0[29]), .Y(n1634) );
  CLKNAND2X2 U1852 ( .A(n1127), .B(n1631), .Y(n1638) );
  XOR2X1 U1853 ( .A(n1639), .B(n1640), .Y(n1127) );
  XOR2X1 U1854 ( .A(n1641), .B(n1642), .Y(n1640) );
  XOR2X1 U1855 ( .A(n1643), .B(C0[28]), .Y(n1639) );
  NAND2BX1 U1856 ( .AN(n1633), .B(n1631), .Y(n1643) );
  XNOR2X1 U1857 ( .A(n1644), .B(n1645), .Y(n1631) );
  XOR2X1 U1858 ( .A(n1646), .B(C0[31]), .Y(n1644) );
  XNOR2X1 U1859 ( .A(n1647), .B(n1648), .Y(n1633) );
  XNOR2X1 U1860 ( .A(C0[30]), .B(n1649), .Y(n1647) );
  OAI221X1 U1861 ( .A0(n1650), .A1(n1257), .B0(n1137), .B1(n1245), .C0(n1651), 
        .Y(Inst_forkAE_L_N33) );
  AOI2BB2X1 U1862 ( .B0(n135), .B1(C1[31]), .A0N(n1247), .A1N(n1134), .Y(n1651) );
  XNOR2X1 U1863 ( .A(n1652), .B(n1653), .Y(n1134) );
  XNOR2X1 U1864 ( .A(n1646), .B(n1654), .Y(n1652) );
  XNOR2X1 U1865 ( .A(Inst_forkAE_CURRENT_KEY_35_), .B(n1655), .Y(n1646) );
  XOR2X1 U1866 ( .A(Inst_forkAE_KEY_INVERSE[82]), .B(
        Inst_forkAE_KEY_INVERSE[147]), .Y(n1655) );
  XOR2X1 U1867 ( .A(n1656), .B(n1657), .Y(n1650) );
  XOR2X1 U1868 ( .A(n712), .B(n1658), .Y(n1657) );
  XOR2X1 U1869 ( .A(Inst_forkAE_KEY_INVERSE[44]), .B(
        Inst_forkAE_KEY_INVERSE[175]), .Y(n1658) );
  XOR2X1 U1870 ( .A(Inst_forkAE_KEY_INVERSE[110]), .B(
        Inst_forkAE_KEY_INVERSE[109]), .Y(n712) );
  XNOR2X1 U1871 ( .A(n1659), .B(n1660), .Y(n1656) );
  XOR2X1 U1872 ( .A(n1661), .B(n837), .Y(n1659) );
  OAI221X1 U1873 ( .A0(n1662), .A1(n1257), .B0(n1663), .B1(n1245), .C0(n1664), 
        .Y(Inst_forkAE_L_N32) );
  AOI22XL U1874 ( .A0(n1138), .A1(n1281), .B0(C1[30]), .B1(n135), .Y(n1664) );
  XNOR2X1 U1875 ( .A(n1665), .B(n1666), .Y(n1138) );
  XOR2X1 U1876 ( .A(n1667), .B(n1649), .Y(n1665) );
  XNOR2X1 U1877 ( .A(n1668), .B(Inst_forkAE_KEY_INVERSE[146]), .Y(n1649) );
  XOR2X1 U1878 ( .A(n355), .B(Inst_forkAE_KEY_INVERSE[81]), .Y(n1668) );
  CLKINVX1 U1879 ( .A(Inst_forkAE_KEY_INVERSE[19]), .Y(n355) );
  XOR2X1 U1880 ( .A(n1669), .B(n1670), .Y(n1662) );
  XOR2X1 U1881 ( .A(n1671), .B(n1672), .Y(n1670) );
  XOR2X1 U1882 ( .A(Inst_forkAE_KEY_INVERSE[174]), .B(
        Inst_forkAE_KEY_INVERSE[109]), .Y(n1672) );
  XOR2X1 U1883 ( .A(Inst_forkAE_KEY_INVERSE[47]), .B(
        Inst_forkAE_KEY_INVERSE[46]), .Y(n1671) );
  XNOR2X1 U1884 ( .A(n1673), .B(n1674), .Y(n1669) );
  XOR2X1 U1885 ( .A(n1675), .B(n837), .Y(n1673) );
  OAI221X1 U1886 ( .A0(n1676), .A1(n1257), .B0(n1145), .B1(n1245), .C0(n1677), 
        .Y(Inst_forkAE_L_N31) );
  AOI2BB2X1 U1887 ( .B0(n135), .B1(C1[29]), .A0N(n1247), .A1N(n1142), .Y(n1677) );
  XOR2X1 U1888 ( .A(n1678), .B(n1679), .Y(n1142) );
  XNOR2X1 U1889 ( .A(C0[34]), .B(n1680), .Y(n1679) );
  NAND2BX1 U1890 ( .AN(C0[33]), .B(n1653), .Y(n1680) );
  XOR2X1 U1891 ( .A(n1681), .B(n1637), .Y(n1678) );
  XNOR2X1 U1892 ( .A(n1682), .B(Inst_forkAE_KEY_INVERSE[145]), .Y(n1637) );
  XOR2X1 U1893 ( .A(n354), .B(Inst_forkAE_KEY_INVERSE[80]), .Y(n1682) );
  CLKINVX1 U1894 ( .A(Inst_forkAE_KEY_INVERSE[18]), .Y(n354) );
  XOR2X1 U1895 ( .A(n1683), .B(n1684), .Y(n1676) );
  XOR2X1 U1896 ( .A(n1685), .B(n1686), .Y(n1684) );
  XOR2X1 U1897 ( .A(n1119), .B(Inst_forkAE_KEY_INVERSE[173]), .Y(n1686) );
  CLKINVX1 U1898 ( .A(C1[34]), .Y(n1119) );
  NAND2BX1 U1899 ( .AN(C1[33]), .B(n1660), .Y(n1685) );
  XOR2X1 U1900 ( .A(n1687), .B(n1688), .Y(n1683) );
  XOR2X1 U1901 ( .A(n466), .B(n837), .Y(n1688) );
  XOR2X1 U1902 ( .A(Inst_forkAE_KEY_INVERSE[108]), .B(
        Inst_forkAE_KEY_INVERSE[111]), .Y(n837) );
  XOR2X1 U1903 ( .A(n554), .B(n549), .Y(n466) );
  CLKINVX1 U1904 ( .A(Inst_forkAE_KEY_INVERSE[46]), .Y(n549) );
  CLKINVX1 U1905 ( .A(Inst_forkAE_KEY_INVERSE[45]), .Y(n554) );
  OAI221X1 U1906 ( .A0(n1689), .A1(n1257), .B0(n1149), .B1(n1245), .C0(n1690), 
        .Y(Inst_forkAE_L_N30) );
  AOI22XL U1907 ( .A0(n1146), .A1(n1281), .B0(n135), .B1(C1[28]), .Y(n1690) );
  XOR2X1 U1908 ( .A(n1691), .B(n1692), .Y(n1146) );
  XNOR2X1 U1909 ( .A(C0[33]), .B(n1693), .Y(n1692) );
  CLKNAND2X2 U1910 ( .A(n1666), .B(n1653), .Y(n1693) );
  XNOR2X1 U1911 ( .A(C0[32]), .B(n1694), .Y(n1653) );
  NOR2X1 U1912 ( .A(C0[34]), .B(C0[35]), .Y(n1694) );
  XNOR2X1 U1913 ( .A(C0[35]), .B(n1695), .Y(n1666) );
  NOR2X1 U1914 ( .A(C0[33]), .B(C0[34]), .Y(n1695) );
  XNOR2X1 U1915 ( .A(n1696), .B(n1642), .Y(n1691) );
  XOR2X1 U1916 ( .A(Inst_forkAE_CURRENT_KEY_96_), .B(n1697), .Y(n1642) );
  XOR2X1 U1917 ( .A(Inst_forkAE_KEY_INVERSE[17]), .B(
        Inst_forkAE_KEY_INVERSE[144]), .Y(n1697) );
  XNOR2X1 U1918 ( .A(n1698), .B(n1541), .Y(n1149) );
  CLKNAND2X2 U1919 ( .A(n1137), .B(n1663), .Y(n1698) );
  XOR2X1 U1920 ( .A(n1699), .B(n1544), .Y(n1137) );
  CLKNAND2X2 U1921 ( .A(n1145), .B(n1663), .Y(n1699) );
  CLKINVX1 U1922 ( .A(n1140), .Y(n1663) );
  XOR2X1 U1923 ( .A(n1700), .B(n1531), .Y(n1140) );
  XOR2X1 U1924 ( .A(C0[37]), .B(C0[5]), .Y(n1531) );
  CLKNAND2X2 U1925 ( .A(n1145), .B(n1541), .Y(n1700) );
  XOR2X1 U1926 ( .A(n1538), .B(n1701), .Y(n1145) );
  NOR2BX1 U1927 ( .AN(n1541), .B(n1544), .Y(n1701) );
  XOR2X1 U1928 ( .A(C0[38]), .B(C0[6]), .Y(n1544) );
  XNOR2X1 U1929 ( .A(C0[39]), .B(C0[7]), .Y(n1541) );
  XNOR2X1 U1930 ( .A(C0[36]), .B(C0[4]), .Y(n1538) );
  XOR2X1 U1931 ( .A(n1702), .B(n1703), .Y(n1689) );
  XOR2X1 U1932 ( .A(n1704), .B(n1705), .Y(n1703) );
  XOR2X1 U1933 ( .A(Inst_forkAE_KEY_INVERSE[172]), .B(
        Inst_forkAE_KEY_INVERSE[111]), .Y(n1705) );
  XOR2X1 U1934 ( .A(Inst_forkAE_KEY_INVERSE[45]), .B(
        Inst_forkAE_KEY_INVERSE[44]), .Y(n1704) );
  XOR2X1 U1935 ( .A(n1706), .B(n1707), .Y(n1702) );
  XNOR2X1 U1936 ( .A(C1[33]), .B(n1708), .Y(n1707) );
  CLKNAND2X2 U1937 ( .A(n1674), .B(n1660), .Y(n1708) );
  XNOR2X1 U1938 ( .A(C1[32]), .B(n1709), .Y(n1660) );
  NOR2X1 U1939 ( .A(C1[35]), .B(C1[34]), .Y(n1709) );
  XNOR2X1 U1940 ( .A(C1[35]), .B(n1710), .Y(n1674) );
  NOR2X1 U1941 ( .A(C1[33]), .B(C1[34]), .Y(n1710) );
  OAI221X1 U1942 ( .A0(n1711), .A1(n1245), .B0(n1151), .B1(n1247), .C0(n1712), 
        .Y(Inst_forkAE_L_N3) );
  AOI22XL U1943 ( .A0(n1249), .A1(n1441), .B0(n135), .B1(C1[1]), .Y(n1712) );
  XOR2X1 U1944 ( .A(n1627), .B(n1713), .Y(n1441) );
  CLKINVX1 U1945 ( .A(n1714), .Y(n1713) );
  XNOR2X1 U1946 ( .A(n1715), .B(n1716), .Y(n1627) );
  XOR2X1 U1947 ( .A(n536), .B(n899), .Y(n1716) );
  XOR2X1 U1948 ( .A(Inst_forkAE_KEY_INVERSE[116]), .B(
        Inst_forkAE_KEY_INVERSE[119]), .Y(n899) );
  XNOR2X1 U1949 ( .A(n501), .B(Inst_forkAE_KEY_INVERSE[54]), .Y(n536) );
  CLKINVX1 U1950 ( .A(Inst_forkAE_KEY_INVERSE[53]), .Y(n501) );
  XOR2X1 U1951 ( .A(n1717), .B(n1718), .Y(n1715) );
  XOR2X1 U1952 ( .A(Inst_forkAE_KEY_INVERSE[181]), .B(C1[50]), .Y(n1718) );
  CLKNAND2X2 U1953 ( .A(n1615), .B(n1044), .Y(n1717) );
  CLKINVX1 U1954 ( .A(C1[49]), .Y(n1044) );
  XOR2X1 U1955 ( .A(n1124), .B(n1719), .Y(n1151) );
  XOR2X1 U1956 ( .A(n1720), .B(n1721), .Y(n1124) );
  XOR2X1 U1957 ( .A(Inst_forkAE_KEY_INVERSE[137]), .B(C0[50]), .Y(n1721) );
  XOR2X1 U1958 ( .A(n1722), .B(n1457), .Y(n1720) );
  XOR2X1 U1959 ( .A(Inst_forkAE_KEY_INVERSE[10]), .B(
        Inst_forkAE_KEY_INVERSE[72]), .Y(n1457) );
  NAND2BX1 U1960 ( .AN(C0[49]), .B(n1617), .Y(n1722) );
  OAI221X1 U1961 ( .A0(n1723), .A1(n1257), .B0(n1157), .B1(n1245), .C0(n1724), 
        .Y(Inst_forkAE_L_N29) );
  AOI22XL U1962 ( .A0(n1154), .A1(n1281), .B0(C1[27]), .B1(n135), .Y(n1724) );
  XOR2X1 U1963 ( .A(n1725), .B(n1726), .Y(n1154) );
  XNOR2X1 U1964 ( .A(n1508), .B(n1727), .Y(n1725) );
  XOR2X1 U1965 ( .A(n334), .B(n1728), .Y(n1508) );
  XOR2X1 U1966 ( .A(Inst_forkAE_KEY_INVERSE[86]), .B(
        Inst_forkAE_KEY_INVERSE[151]), .Y(n1728) );
  CLKINVX1 U1967 ( .A(Inst_forkAE_CURRENT_KEY_47_), .Y(n334) );
  XOR2X1 U1968 ( .A(n1729), .B(n1730), .Y(n1723) );
  XOR2X1 U1969 ( .A(n908), .B(n1731), .Y(n1730) );
  XOR2X1 U1970 ( .A(Inst_forkAE_KEY_INVERSE[32]), .B(
        Inst_forkAE_KEY_INVERSE[163]), .Y(n1731) );
  XOR2X1 U1971 ( .A(Inst_forkAE_KEY_INVERSE[98]), .B(
        Inst_forkAE_KEY_INVERSE[97]), .Y(n908) );
  XOR2X1 U1972 ( .A(n1732), .B(n1733), .Y(n1729) );
  XOR2X1 U1973 ( .A(n1734), .B(n919), .Y(n1732) );
  OAI221X1 U1974 ( .A0(n1257), .A1(n1735), .B0(n1162), .B1(n1245), .C0(n1736), 
        .Y(Inst_forkAE_L_N28) );
  AOI2BB2X1 U1975 ( .B0(n135), .B1(C1[26]), .A0N(n1247), .A1N(n1159), .Y(n1736) );
  XNOR2X1 U1976 ( .A(n1737), .B(n1738), .Y(n1159) );
  XNOR2X1 U1977 ( .A(n1739), .B(n1740), .Y(n1738) );
  XOR2X1 U1978 ( .A(n181), .B(Inst_forkAE_KEY_INVERSE[150]), .Y(n1740) );
  XNOR2X1 U1979 ( .A(n1741), .B(n1512), .Y(n1737) );
  XOR2X1 U1980 ( .A(Inst_forkAE_KEY_INVERSE[23]), .B(
        Inst_forkAE_KEY_INVERSE[85]), .Y(n1512) );
  XOR2X1 U1981 ( .A(n1742), .B(n1743), .Y(n1735) );
  XNOR2X1 U1982 ( .A(n1744), .B(n1745), .Y(n1743) );
  XOR2X1 U1983 ( .A(n1746), .B(n1747), .Y(n1744) );
  XOR2X1 U1984 ( .A(Inst_forkAE_KEY_INVERSE[35]), .B(n1748), .Y(n1747) );
  XOR2X1 U1985 ( .A(n180), .B(Inst_forkAE_KEY_INVERSE[97]), .Y(n1748) );
  XOR2X1 U1986 ( .A(n1749), .B(n1750), .Y(n1746) );
  XNOR2X1 U1987 ( .A(n1751), .B(Inst_forkAE_KEY_INVERSE[34]), .Y(n1749) );
  XNOR2X1 U1988 ( .A(n919), .B(Inst_forkAE_KEY_INVERSE[162]), .Y(n1742) );
  OAI221X1 U1989 ( .A0(n1752), .A1(n1257), .B0(n1166), .B1(n1245), .C0(n1753), 
        .Y(Inst_forkAE_L_N27) );
  AOI22XL U1990 ( .A0(n1163), .A1(n1281), .B0(C1[25]), .B1(n135), .Y(n1753) );
  XOR2X1 U1991 ( .A(n1754), .B(n1755), .Y(n1163) );
  XOR2X1 U1992 ( .A(C0[46]), .B(n1756), .Y(n1755) );
  XOR2X1 U1993 ( .A(Inst_forkAE_KEY_INVERSE[149]), .B(Inst_forkAE_CONST_ENC_5_), .Y(n1756) );
  XOR2X1 U1994 ( .A(n1757), .B(n1497), .Y(n1754) );
  XOR2X1 U1995 ( .A(Inst_forkAE_KEY_INVERSE[22]), .B(
        Inst_forkAE_KEY_INVERSE[84]), .Y(n1497) );
  XNOR2X1 U1996 ( .A(n1758), .B(n1759), .Y(n1757) );
  NOR2X1 U1997 ( .A(C0[45]), .B(n1726), .Y(n1759) );
  XOR2X1 U1998 ( .A(n1760), .B(n1761), .Y(n1752) );
  XOR2X1 U1999 ( .A(n1762), .B(n1763), .Y(n1761) );
  XOR2X1 U2000 ( .A(n1764), .B(n561), .Y(n1763) );
  XOR2X1 U2001 ( .A(n460), .B(Inst_forkAE_KEY_INVERSE[34]), .Y(n561) );
  CLKINVX1 U2002 ( .A(Inst_forkAE_KEY_INVERSE[33]), .Y(n460) );
  NAND2BX1 U2003 ( .AN(C1[45]), .B(n1765), .Y(n1764) );
  XOR2X1 U2004 ( .A(Inst_forkAE_KEY_INVERSE[161]), .B(C1[46]), .Y(n1762) );
  XOR2X1 U2005 ( .A(n1766), .B(n1767), .Y(n1760) );
  XNOR2X1 U2006 ( .A(n919), .B(n1768), .Y(n1767) );
  XOR2X1 U2007 ( .A(n891), .B(n709), .Y(n919) );
  CLKINVX1 U2008 ( .A(Inst_forkAE_KEY_INVERSE[99]), .Y(n709) );
  CLKINVX1 U2009 ( .A(Inst_forkAE_KEY_INVERSE[96]), .Y(n891) );
  XOR2X1 U2010 ( .A(n1769), .B(n1751), .Y(n1766) );
  XNOR2X1 U2011 ( .A(n132), .B(n1770), .Y(n1751) );
  OAI221X1 U2012 ( .A0(n1257), .A1(n1771), .B0(n1170), .B1(n1245), .C0(n1772), 
        .Y(Inst_forkAE_L_N26) );
  AOI22XL U2013 ( .A0(n1281), .A1(n1167), .B0(C1[24]), .B1(n135), .Y(n1772) );
  XNOR2X1 U2014 ( .A(n1773), .B(n1774), .Y(n1167) );
  XOR2X1 U2015 ( .A(C0[45]), .B(n1775), .Y(n1774) );
  XOR2X1 U2016 ( .A(n180), .B(Inst_forkAE_KEY_INVERSE[148]), .Y(n1775) );
  XOR2X1 U2017 ( .A(n1776), .B(n1505), .Y(n1773) );
  XOR2X1 U2018 ( .A(Inst_forkAE_CURRENT_KEY_108_), .B(
        Inst_forkAE_KEY_INVERSE[21]), .Y(n1505) );
  XOR2X1 U2019 ( .A(n1777), .B(n1778), .Y(n1776) );
  NOR2X1 U2020 ( .A(n1726), .B(n1741), .Y(n1778) );
  XNOR2X1 U2021 ( .A(n1302), .B(n1779), .Y(n1741) );
  NOR2X1 U2022 ( .A(C0[45]), .B(C0[46]), .Y(n1779) );
  CLKINVX1 U2023 ( .A(C0[47]), .Y(n1302) );
  XOR2X1 U2024 ( .A(C0[44]), .B(n1780), .Y(n1726) );
  NOR2X1 U2025 ( .A(C0[46]), .B(C0[47]), .Y(n1780) );
  XNOR2X1 U2026 ( .A(n1781), .B(n1605), .Y(n1170) );
  CLKNAND2X2 U2027 ( .A(n1157), .B(n1162), .Y(n1781) );
  XOR2X1 U2028 ( .A(n1782), .B(n1608), .Y(n1157) );
  CLKNAND2X2 U2029 ( .A(n1162), .B(n1166), .Y(n1782) );
  XOR2X1 U2030 ( .A(n1783), .B(n1596), .Y(n1162) );
  XOR2X1 U2031 ( .A(C0[1]), .B(C0[33]), .Y(n1596) );
  CLKNAND2X2 U2032 ( .A(n1166), .B(n1605), .Y(n1783) );
  XNOR2X1 U2033 ( .A(n1601), .B(n1784), .Y(n1166) );
  NOR2BX1 U2034 ( .AN(n1605), .B(n1608), .Y(n1784) );
  XOR2X1 U2035 ( .A(C0[2]), .B(C0[34]), .Y(n1608) );
  XNOR2X1 U2036 ( .A(C0[35]), .B(C0[3]), .Y(n1605) );
  XOR2X1 U2037 ( .A(C0[0]), .B(C0[32]), .Y(n1601) );
  XOR2X1 U2038 ( .A(n1785), .B(n1786), .Y(n1771) );
  XOR2X1 U2039 ( .A(C1[45]), .B(n431), .Y(n1786) );
  CLKINVX1 U2040 ( .A(Inst_forkAE_KEY_INVERSE[32]), .Y(n431) );
  XOR2X1 U2041 ( .A(n1787), .B(n1788), .Y(n1785) );
  XOR2X1 U2042 ( .A(n1789), .B(n1790), .Y(n1788) );
  XOR2X1 U2043 ( .A(Inst_forkAE_KEY_INVERSE[160]), .B(Inst_forkAE_CONST_ENC_5_), .Y(n1790) );
  XOR2X1 U2044 ( .A(Inst_forkAE_KEY_INVERSE[99]), .B(
        Inst_forkAE_KEY_INVERSE[33]), .Y(n1789) );
  XOR2X1 U2045 ( .A(n1791), .B(n1792), .Y(n1787) );
  XOR2X1 U2046 ( .A(n1793), .B(n1794), .Y(n1792) );
  NOR2X1 U2047 ( .A(n1733), .B(n1750), .Y(n1793) );
  XOR2X1 U2048 ( .A(C1[47]), .B(n1795), .Y(n1750) );
  NOR2X1 U2049 ( .A(C1[45]), .B(C1[46]), .Y(n1795) );
  CLKINVX1 U2050 ( .A(n1765), .Y(n1733) );
  XNOR2X1 U2051 ( .A(C1[44]), .B(n1796), .Y(n1765) );
  NOR2X1 U2052 ( .A(C1[46]), .B(C1[47]), .Y(n1796) );
  XOR2X1 U2053 ( .A(n1797), .B(n1770), .Y(n1791) );
  XOR2X1 U2054 ( .A(Inst_forkAE_CONST_ENC_1_), .B(Inst_forkAE_CONST_ENC_2_), 
        .Y(n1770) );
  OAI221X1 U2055 ( .A0(n1798), .A1(n1257), .B0(n1175), .B1(n1245), .C0(n1799), 
        .Y(Inst_forkAE_L_N25) );
  AOI2BB2X1 U2056 ( .B0(n135), .B1(C1[23]), .A0N(n1247), .A1N(n1172), .Y(n1799) );
  XNOR2X1 U2057 ( .A(n1800), .B(n1801), .Y(n1172) );
  XNOR2X1 U2058 ( .A(n1542), .B(n1371), .Y(n1800) );
  XNOR2X1 U2059 ( .A(Inst_forkAE_CURRENT_KEY_43_), .B(n1802), .Y(n1542) );
  XOR2X1 U2060 ( .A(Inst_forkAE_KEY_INVERSE[70]), .B(
        Inst_forkAE_KEY_INVERSE[135]), .Y(n1802) );
  XOR2X1 U2061 ( .A(n1803), .B(n1804), .Y(n1798) );
  XOR2X1 U2062 ( .A(Inst_forkAE_KEY_INVERSE[126]), .B(n1805), .Y(n1804) );
  XOR2X1 U2063 ( .A(Inst_forkAE_KEY_INVERSE[60]), .B(
        Inst_forkAE_KEY_INVERSE[191]), .Y(n1805) );
  XOR2X1 U2064 ( .A(n1806), .B(n1807), .Y(n1803) );
  XNOR2X1 U2065 ( .A(n1374), .B(n1808), .Y(n1806) );
  OAI221X1 U2066 ( .A0(n1809), .A1(n1257), .B0(n1179), .B1(n1245), .C0(n1810), 
        .Y(Inst_forkAE_L_N24) );
  AOI22XL U2067 ( .A0(n1176), .A1(n1281), .B0(C1[22]), .B1(n135), .Y(n1810) );
  XNOR2X1 U2068 ( .A(n1811), .B(n1812), .Y(n1176) );
  XOR2X1 U2069 ( .A(n1380), .B(n1545), .Y(n1811) );
  XNOR2X1 U2070 ( .A(n1813), .B(Inst_forkAE_KEY_INVERSE[134]), .Y(n1545) );
  XOR2X1 U2071 ( .A(n601), .B(Inst_forkAE_KEY_INVERSE[7]), .Y(n1813) );
  CLKINVX1 U2072 ( .A(Inst_forkAE_KEY_INVERSE[69]), .Y(n601) );
  XOR2X1 U2073 ( .A(n1814), .B(n1815), .Y(n1809) );
  XOR2X1 U2074 ( .A(Inst_forkAE_KEY_INVERSE[190]), .B(n1816), .Y(n1815) );
  XOR2X1 U2075 ( .A(Inst_forkAE_KEY_INVERSE[63]), .B(
        Inst_forkAE_KEY_INVERSE[62]), .Y(n1816) );
  XNOR2X1 U2076 ( .A(n1817), .B(n1818), .Y(n1814) );
  XOR2X1 U2077 ( .A(n1807), .B(n1384), .Y(n1817) );
  XNOR2X1 U2078 ( .A(n619), .B(n940), .Y(n1807) );
  CLKINVX1 U2079 ( .A(Inst_forkAE_KEY_INVERSE[125]), .Y(n619) );
  OAI221X1 U2080 ( .A0(n1257), .A1(n1819), .B0(n1183), .B1(n1245), .C0(n1820), 
        .Y(Inst_forkAE_L_N23) );
  AOI22XL U2081 ( .A0(n1281), .A1(n1180), .B0(C1[21]), .B1(n135), .Y(n1820) );
  XNOR2X1 U2082 ( .A(n1821), .B(n1822), .Y(n1180) );
  XOR2X1 U2083 ( .A(n1823), .B(n1824), .Y(n1822) );
  XNOR2X1 U2084 ( .A(Inst_forkAE_KEY_INVERSE[133]), .B(C0[42]), .Y(n1824) );
  NAND2BX1 U2085 ( .AN(C0[41]), .B(n1801), .Y(n1823) );
  XNOR2X1 U2086 ( .A(n1390), .B(n1530), .Y(n1821) );
  XOR2X1 U2087 ( .A(Inst_forkAE_KEY_INVERSE[68]), .B(
        Inst_forkAE_KEY_INVERSE[6]), .Y(n1530) );
  XNOR2X1 U2088 ( .A(n1825), .B(C0[30]), .Y(n1390) );
  NAND2BX1 U2089 ( .AN(C0[29]), .B(n1371), .Y(n1825) );
  XOR2X1 U2090 ( .A(n1826), .B(n1827), .Y(n1819) );
  XOR2X1 U2091 ( .A(n1395), .B(n1828), .Y(n1827) );
  XNOR2X1 U2092 ( .A(n940), .B(n584), .Y(n1828) );
  XNOR2X1 U2093 ( .A(n448), .B(Inst_forkAE_KEY_INVERSE[62]), .Y(n584) );
  CLKINVX1 U2094 ( .A(Inst_forkAE_KEY_INVERSE[61]), .Y(n448) );
  XNOR2X1 U2095 ( .A(n829), .B(Inst_forkAE_KEY_INVERSE[127]), .Y(n940) );
  CLKINVX1 U2096 ( .A(Inst_forkAE_KEY_INVERSE[124]), .Y(n829) );
  XOR2X1 U2097 ( .A(n1829), .B(C1[30]), .Y(n1395) );
  CLKNAND2X2 U2098 ( .A(n1374), .B(n1141), .Y(n1829) );
  CLKINVX1 U2099 ( .A(C1[29]), .Y(n1141) );
  XOR2X1 U2100 ( .A(n1830), .B(n1831), .Y(n1826) );
  XNOR2X1 U2101 ( .A(C1[42]), .B(Inst_forkAE_KEY_INVERSE[189]), .Y(n1831) );
  NAND2BX1 U2102 ( .AN(C1[41]), .B(n1808), .Y(n1830) );
  OAI221X1 U2103 ( .A0(n1832), .A1(n1257), .B0(n1187), .B1(n1245), .C0(n1833), 
        .Y(Inst_forkAE_L_N22) );
  AOI22XL U2104 ( .A0(n1184), .A1(n1281), .B0(C1[20]), .B1(n135), .Y(n1833) );
  XOR2X1 U2105 ( .A(n1834), .B(n1835), .Y(n1184) );
  XNOR2X1 U2106 ( .A(C0[41]), .B(n1836), .Y(n1835) );
  CLKNAND2X2 U2107 ( .A(n1812), .B(n1801), .Y(n1836) );
  XNOR2X1 U2108 ( .A(C0[40]), .B(n1837), .Y(n1801) );
  NOR2X1 U2109 ( .A(C0[42]), .B(C0[43]), .Y(n1837) );
  XNOR2X1 U2110 ( .A(C0[43]), .B(n1838), .Y(n1812) );
  NOR2X1 U2111 ( .A(C0[41]), .B(C0[42]), .Y(n1838) );
  XNOR2X1 U2112 ( .A(n1402), .B(n1537), .Y(n1834) );
  XOR2X1 U2113 ( .A(Inst_forkAE_CURRENT_KEY_104_), .B(n1839), .Y(n1537) );
  XOR2X1 U2114 ( .A(Inst_forkAE_KEY_INVERSE[5]), .B(
        Inst_forkAE_KEY_INVERSE[132]), .Y(n1839) );
  XNOR2X1 U2115 ( .A(n1840), .B(C0[29]), .Y(n1402) );
  CLKNAND2X2 U2116 ( .A(n1380), .B(n1371), .Y(n1840) );
  XNOR2X1 U2117 ( .A(C0[28]), .B(n1841), .Y(n1371) );
  NOR2X1 U2118 ( .A(C0[30]), .B(C0[31]), .Y(n1841) );
  XNOR2X1 U2119 ( .A(C0[31]), .B(n1842), .Y(n1380) );
  NOR2X1 U2120 ( .A(C0[29]), .B(C0[30]), .Y(n1842) );
  XOR2X1 U2121 ( .A(n1843), .B(n1844), .Y(n1187) );
  CLKNAND2X2 U2122 ( .A(n1175), .B(n1179), .Y(n1843) );
  XOR2X1 U2123 ( .A(n1845), .B(n1648), .Y(n1175) );
  CLKNAND2X2 U2124 ( .A(n1179), .B(n1183), .Y(n1845) );
  XOR2X1 U2125 ( .A(n1846), .B(n1636), .Y(n1179) );
  XOR2X1 U2126 ( .A(C0[13]), .B(C0[45]), .Y(n1636) );
  CLKNAND2X2 U2127 ( .A(n1183), .B(n1645), .Y(n1846) );
  CLKINVX1 U2128 ( .A(n1844), .Y(n1645) );
  XNOR2X1 U2129 ( .A(n1641), .B(n1847), .Y(n1183) );
  NOR2X1 U2130 ( .A(n1648), .B(n1844), .Y(n1847) );
  XOR2X1 U2131 ( .A(C0[15]), .B(C0[47]), .Y(n1844) );
  XOR2X1 U2132 ( .A(C0[14]), .B(C0[46]), .Y(n1648) );
  XOR2X1 U2133 ( .A(C0[12]), .B(C0[44]), .Y(n1641) );
  XOR2X1 U2134 ( .A(n1848), .B(n1849), .Y(n1832) );
  XOR2X1 U2135 ( .A(n1850), .B(n1851), .Y(n1849) );
  XOR2X1 U2136 ( .A(Inst_forkAE_KEY_INVERSE[188]), .B(
        Inst_forkAE_KEY_INVERSE[127]), .Y(n1851) );
  XOR2X1 U2137 ( .A(Inst_forkAE_KEY_INVERSE[61]), .B(
        Inst_forkAE_KEY_INVERSE[60]), .Y(n1850) );
  XOR2X1 U2138 ( .A(n1425), .B(n1852), .Y(n1848) );
  XNOR2X1 U2139 ( .A(C1[41]), .B(n1853), .Y(n1852) );
  CLKNAND2X2 U2140 ( .A(n1818), .B(n1808), .Y(n1853) );
  XOR2X1 U2141 ( .A(n1088), .B(n1854), .Y(n1808) );
  NOR2X1 U2142 ( .A(C1[42]), .B(C1[43]), .Y(n1854) );
  CLKINVX1 U2143 ( .A(C1[40]), .Y(n1088) );
  XNOR2X1 U2144 ( .A(C1[43]), .B(n1855), .Y(n1818) );
  NOR2X1 U2145 ( .A(C1[41]), .B(C1[42]), .Y(n1855) );
  XOR2X1 U2146 ( .A(n1856), .B(C1[29]), .Y(n1425) );
  CLKNAND2X2 U2147 ( .A(n1384), .B(n1374), .Y(n1856) );
  XNOR2X1 U2148 ( .A(C1[28]), .B(n1857), .Y(n1374) );
  NOR2X1 U2149 ( .A(C1[30]), .B(C1[31]), .Y(n1857) );
  XOR2X1 U2150 ( .A(n1133), .B(n1858), .Y(n1384) );
  NOR2X1 U2151 ( .A(C1[30]), .B(C1[29]), .Y(n1858) );
  CLKINVX1 U2152 ( .A(C1[31]), .Y(n1133) );
  OAI221X1 U2153 ( .A0(n1859), .A1(n1257), .B0(n1191), .B1(n1245), .C0(n1860), 
        .Y(Inst_forkAE_L_N21) );
  AOI22XL U2154 ( .A0(n1188), .A1(n1281), .B0(C1[19]), .B1(n135), .Y(n1860) );
  XNOR2X1 U2155 ( .A(n1861), .B(n1862), .Y(n1188) );
  XNOR2X1 U2156 ( .A(n1606), .B(n1475), .Y(n1861) );
  XNOR2X1 U2157 ( .A(Inst_forkAE_CURRENT_KEY_39_), .B(n1863), .Y(n1606) );
  XOR2X1 U2158 ( .A(Inst_forkAE_KEY_INVERSE[78]), .B(
        Inst_forkAE_KEY_INVERSE[143]), .Y(n1863) );
  XOR2X1 U2159 ( .A(n1864), .B(n1865), .Y(n1859) );
  XOR2X1 U2160 ( .A(Inst_forkAE_KEY_INVERSE[122]), .B(n1866), .Y(n1865) );
  XOR2X1 U2161 ( .A(Inst_forkAE_KEY_INVERSE[56]), .B(
        Inst_forkAE_KEY_INVERSE[187]), .Y(n1866) );
  XOR2X1 U2162 ( .A(n1867), .B(n1868), .Y(n1864) );
  CLKINVX1 U2163 ( .A(n1869), .Y(n1868) );
  XNOR2X1 U2164 ( .A(n1473), .B(n1870), .Y(n1867) );
  OAI221X1 U2165 ( .A0(n1871), .A1(n1257), .B0(n1195), .B1(n1245), .C0(n1872), 
        .Y(Inst_forkAE_L_N20) );
  AOI22XL U2166 ( .A0(n1192), .A1(n1281), .B0(C1[18]), .B1(n135), .Y(n1872) );
  XNOR2X1 U2167 ( .A(n1873), .B(n1874), .Y(n1192) );
  XOR2X1 U2168 ( .A(n1567), .B(n1609), .Y(n1873) );
  XNOR2X1 U2169 ( .A(n1875), .B(Inst_forkAE_KEY_INVERSE[142]), .Y(n1609) );
  XOR2X1 U2170 ( .A(n268), .B(Inst_forkAE_KEY_INVERSE[77]), .Y(n1875) );
  CLKINVX1 U2171 ( .A(Inst_forkAE_KEY_INVERSE[15]), .Y(n268) );
  XOR2X1 U2172 ( .A(n1876), .B(n1877), .Y(n1871) );
  XOR2X1 U2173 ( .A(Inst_forkAE_KEY_INVERSE[186]), .B(n1878), .Y(n1877) );
  XOR2X1 U2174 ( .A(Inst_forkAE_KEY_INVERSE[59]), .B(
        Inst_forkAE_KEY_INVERSE[58]), .Y(n1878) );
  XNOR2X1 U2175 ( .A(n1879), .B(n1880), .Y(n1876) );
  XOR2X1 U2176 ( .A(n1869), .B(n1565), .Y(n1879) );
  CLKINVX1 U2177 ( .A(n1881), .Y(n1565) );
  XOR2X1 U2178 ( .A(n647), .B(n607), .Y(n1869) );
  CLKINVX1 U2179 ( .A(Inst_forkAE_KEY_INVERSE[121]), .Y(n647) );
  OAI221X1 U2180 ( .A0(n1199), .A1(n1245), .B0(n1882), .B1(n1247), .C0(n1883), 
        .Y(Inst_forkAE_L_N2) );
  AOI22XL U2181 ( .A0(n1249), .A1(n1466), .B0(C1[0]), .B1(n135), .Y(n1883) );
  XOR2X1 U2182 ( .A(n1629), .B(n1884), .Y(n1466) );
  CLKINVX1 U2183 ( .A(n1885), .Y(n1884) );
  XNOR2X1 U2184 ( .A(n1886), .B(n1887), .Y(n1629) );
  XOR2X1 U2185 ( .A(Inst_forkAE_KEY_INVERSE[180]), .B(n1888), .Y(n1887) );
  XOR2X1 U2186 ( .A(Inst_forkAE_KEY_INVERSE[53]), .B(
        Inst_forkAE_KEY_INVERSE[52]), .Y(n1888) );
  XOR2X1 U2187 ( .A(n1889), .B(n1890), .Y(n1886) );
  XOR2X1 U2188 ( .A(Inst_forkAE_KEY_INVERSE[119]), .B(C1[49]), .Y(n1890) );
  CLKNAND2X2 U2189 ( .A(n1622), .B(n1615), .Y(n1889) );
  XNOR2X1 U2190 ( .A(C1[48]), .B(n1891), .Y(n1615) );
  NOR2X1 U2191 ( .A(C1[51]), .B(C1[50]), .Y(n1891) );
  XNOR2X1 U2192 ( .A(C1[51]), .B(n1892), .Y(n1622) );
  NOR2X1 U2193 ( .A(C1[49]), .B(C1[50]), .Y(n1892) );
  CLKINVX1 U2194 ( .A(n1196), .Y(n1882) );
  XOR2X1 U2195 ( .A(n1129), .B(n1893), .Y(n1196) );
  CLKINVX1 U2196 ( .A(n1894), .Y(n1893) );
  XOR2X1 U2197 ( .A(n1895), .B(n1896), .Y(n1129) );
  XOR2X1 U2198 ( .A(Inst_forkAE_KEY_INVERSE[136]), .B(C0[49]), .Y(n1896) );
  XOR2X1 U2199 ( .A(n1897), .B(n1461), .Y(n1895) );
  XOR2X1 U2200 ( .A(Inst_forkAE_CURRENT_KEY_112_), .B(
        Inst_forkAE_KEY_INVERSE[9]), .Y(n1461) );
  CLKNAND2X2 U2201 ( .A(n1624), .B(n1617), .Y(n1897) );
  XNOR2X1 U2202 ( .A(C0[48]), .B(n1898), .Y(n1617) );
  NOR2X1 U2203 ( .A(C0[50]), .B(C0[51]), .Y(n1898) );
  XNOR2X1 U2204 ( .A(C0[51]), .B(n1899), .Y(n1624) );
  NOR2X1 U2205 ( .A(C0[49]), .B(C0[50]), .Y(n1899) );
  XOR2X1 U2206 ( .A(n1900), .B(n1901), .Y(n1199) );
  CLKNAND2X2 U2207 ( .A(n1057), .B(n1105), .Y(n1900) );
  XOR2X1 U2208 ( .A(n1902), .B(n1903), .Y(n1057) );
  CLKNAND2X2 U2209 ( .A(n1105), .B(n1711), .Y(n1902) );
  XOR2X1 U2210 ( .A(n1904), .B(n1905), .Y(n1105) );
  XOR2X1 U2211 ( .A(C0[5]), .B(C0[53]), .Y(n1905) );
  OR2X1 U2212 ( .A(n1901), .B(n1153), .Y(n1904) );
  CLKINVX1 U2213 ( .A(n1711), .Y(n1153) );
  XOR2X1 U2214 ( .A(n1906), .B(n1907), .Y(n1711) );
  NOR2X1 U2215 ( .A(n1901), .B(n1903), .Y(n1907) );
  XOR2X1 U2216 ( .A(C0[54]), .B(C0[6]), .Y(n1903) );
  XNOR2X1 U2217 ( .A(C0[4]), .B(C0[52]), .Y(n1906) );
  XOR2X1 U2218 ( .A(C0[55]), .B(C0[7]), .Y(n1901) );
  OAI221X1 U2219 ( .A0(n1908), .A1(n1257), .B0(n1203), .B1(n1245), .C0(n1909), 
        .Y(Inst_forkAE_L_N19) );
  AOI22XL U2220 ( .A0(n1200), .A1(n1281), .B0(C1[17]), .B1(n135), .Y(n1909) );
  XOR2X1 U2221 ( .A(n1910), .B(n1911), .Y(n1200) );
  XOR2X1 U2222 ( .A(n1418), .B(n1912), .Y(n1911) );
  NAND2BX1 U2223 ( .AN(C0[37]), .B(n1862), .Y(n1912) );
  CLKINVX1 U2224 ( .A(C0[38]), .Y(n1418) );
  XNOR2X1 U2225 ( .A(n1719), .B(n1597), .Y(n1910) );
  XNOR2X1 U2226 ( .A(n1913), .B(Inst_forkAE_KEY_INVERSE[141]), .Y(n1597) );
  XOR2X1 U2227 ( .A(n267), .B(Inst_forkAE_KEY_INVERSE[76]), .Y(n1913) );
  CLKINVX1 U2228 ( .A(Inst_forkAE_KEY_INVERSE[14]), .Y(n267) );
  XNOR2X1 U2229 ( .A(n1914), .B(C0[26]), .Y(n1719) );
  NAND2BX1 U2230 ( .AN(C0[25]), .B(n1475), .Y(n1914) );
  XOR2X1 U2231 ( .A(n1915), .B(n1916), .Y(n1908) );
  XOR2X1 U2232 ( .A(n1917), .B(n1918), .Y(n1916) );
  XNOR2X1 U2233 ( .A(C1[38]), .B(Inst_forkAE_KEY_INVERSE[185]), .Y(n1918) );
  CLKNAND2X2 U2234 ( .A(n1870), .B(n1106), .Y(n1917) );
  XOR2X1 U2235 ( .A(n1714), .B(n1919), .Y(n1915) );
  XOR2X1 U2236 ( .A(n211), .B(n607), .Y(n1919) );
  XOR2X1 U2237 ( .A(Inst_forkAE_KEY_INVERSE[120]), .B(
        Inst_forkAE_KEY_INVERSE[123]), .Y(n607) );
  XOR2X1 U2238 ( .A(n479), .B(n474), .Y(n211) );
  CLKINVX1 U2239 ( .A(Inst_forkAE_KEY_INVERSE[58]), .Y(n474) );
  CLKINVX1 U2240 ( .A(Inst_forkAE_KEY_INVERSE[57]), .Y(n479) );
  XOR2X1 U2241 ( .A(n1920), .B(C1[26]), .Y(n1714) );
  NAND2BX1 U2242 ( .AN(C1[25]), .B(n1473), .Y(n1920) );
  OAI221X1 U2243 ( .A0(n1921), .A1(n1257), .B0(n1207), .B1(n1245), .C0(n1922), 
        .Y(Inst_forkAE_L_N18) );
  AOI22XL U2244 ( .A0(n1204), .A1(n1281), .B0(C1[16]), .B1(n135), .Y(n1922) );
  CLKINVX1 U2245 ( .A(n1247), .Y(n1281) );
  XOR2X1 U2246 ( .A(n1923), .B(n1924), .Y(n1204) );
  XNOR2X1 U2247 ( .A(C0[37]), .B(n1925), .Y(n1924) );
  CLKNAND2X2 U2248 ( .A(n1874), .B(n1862), .Y(n1925) );
  XNOR2X1 U2249 ( .A(C0[36]), .B(n1926), .Y(n1862) );
  NOR2X1 U2250 ( .A(C0[38]), .B(C0[39]), .Y(n1926) );
  XNOR2X1 U2251 ( .A(C0[39]), .B(n1927), .Y(n1874) );
  NOR2X1 U2252 ( .A(C0[37]), .B(C0[38]), .Y(n1927) );
  XOR2X1 U2253 ( .A(n1894), .B(n1602), .Y(n1923) );
  XOR2X1 U2254 ( .A(Inst_forkAE_CURRENT_KEY_100_), .B(n1928), .Y(n1602) );
  XOR2X1 U2255 ( .A(Inst_forkAE_KEY_INVERSE[140]), .B(
        Inst_forkAE_KEY_INVERSE[13]), .Y(n1928) );
  XOR2X1 U2256 ( .A(n1929), .B(C0[25]), .Y(n1894) );
  CLKNAND2X2 U2257 ( .A(n1567), .B(n1475), .Y(n1929) );
  XNOR2X1 U2258 ( .A(C0[24]), .B(n1930), .Y(n1475) );
  NOR2X1 U2259 ( .A(C0[26]), .B(C0[27]), .Y(n1930) );
  XNOR2X1 U2260 ( .A(C0[27]), .B(n1931), .Y(n1567) );
  NOR2X1 U2261 ( .A(C0[25]), .B(C0[26]), .Y(n1931) );
  XOR2X1 U2262 ( .A(n1932), .B(n1933), .Y(n1207) );
  CLKNAND2X2 U2263 ( .A(n1191), .B(n1195), .Y(n1932) );
  XOR2X1 U2264 ( .A(n1934), .B(n1511), .Y(n1191) );
  CLKNAND2X2 U2265 ( .A(n1195), .B(n1203), .Y(n1934) );
  XOR2X1 U2266 ( .A(n1935), .B(n1495), .Y(n1195) );
  XOR2X1 U2267 ( .A(C0[41]), .B(C0[9]), .Y(n1495) );
  CLKNAND2X2 U2268 ( .A(n1203), .B(n1507), .Y(n1935) );
  CLKINVX1 U2269 ( .A(n1933), .Y(n1507) );
  XOR2X1 U2270 ( .A(n1503), .B(n1936), .Y(n1203) );
  NOR2X1 U2271 ( .A(n1511), .B(n1933), .Y(n1936) );
  XOR2X1 U2272 ( .A(C0[11]), .B(C0[43]), .Y(n1933) );
  XOR2X1 U2273 ( .A(C0[10]), .B(C0[42]), .Y(n1511) );
  XNOR2X1 U2274 ( .A(C0[40]), .B(C0[8]), .Y(n1503) );
  XOR2X1 U2275 ( .A(n1937), .B(n1938), .Y(n1921) );
  XOR2X1 U2276 ( .A(n1939), .B(n1940), .Y(n1938) );
  XOR2X1 U2277 ( .A(Inst_forkAE_KEY_INVERSE[184]), .B(
        Inst_forkAE_KEY_INVERSE[123]), .Y(n1940) );
  XOR2X1 U2278 ( .A(Inst_forkAE_KEY_INVERSE[57]), .B(
        Inst_forkAE_KEY_INVERSE[56]), .Y(n1939) );
  XOR2X1 U2279 ( .A(n1885), .B(n1941), .Y(n1937) );
  XOR2X1 U2280 ( .A(n1106), .B(n1942), .Y(n1941) );
  CLKNAND2X2 U2281 ( .A(n1880), .B(n1870), .Y(n1942) );
  XNOR2X1 U2282 ( .A(C1[36]), .B(n1943), .Y(n1870) );
  NOR2X1 U2283 ( .A(C1[38]), .B(C1[39]), .Y(n1943) );
  XNOR2X1 U2284 ( .A(C1[39]), .B(n1944), .Y(n1880) );
  NOR2X1 U2285 ( .A(C1[38]), .B(C1[37]), .Y(n1944) );
  CLKINVX1 U2286 ( .A(C1[37]), .Y(n1106) );
  XOR2X1 U2287 ( .A(n1945), .B(C1[25]), .Y(n1885) );
  CLKNAND2X2 U2288 ( .A(n1881), .B(n1473), .Y(n1945) );
  XNOR2X1 U2289 ( .A(C1[24]), .B(n1946), .Y(n1473) );
  NOR2X1 U2290 ( .A(C1[27]), .B(C1[26]), .Y(n1946) );
  XNOR2X1 U2291 ( .A(C1[27]), .B(n1947), .Y(n1881) );
  NOR2X1 U2292 ( .A(C1[25]), .B(C1[26]), .Y(n1947) );
  OAI221X1 U2293 ( .A0(n1211), .A1(n1245), .B0(n1212), .B1(n1247), .C0(n1948), 
        .Y(Inst_forkAE_L_N17) );
  AOI2BB2X1 U2294 ( .B0(C1[15]), .B1(n135), .A0N(n1263), .A1N(n1257), .Y(n1948) );
  XNOR2X1 U2295 ( .A(n1477), .B(n1949), .Y(n1263) );
  XOR2X1 U2296 ( .A(n1950), .B(n1951), .Y(n1477) );
  XOR2X1 U2297 ( .A(n1952), .B(n1953), .Y(n1951) );
  XOR2X1 U2298 ( .A(Inst_forkAE_KEY_INVERSE[171]), .B(Inst_forkAE_CONST_ENC_1_), .Y(n1953) );
  XOR2X1 U2299 ( .A(n180), .B(Inst_forkAE_KEY_INVERSE[40]), .Y(n1952) );
  XOR2X1 U2300 ( .A(n1954), .B(n1955), .Y(n1950) );
  XOR2X1 U2301 ( .A(n816), .B(n827), .Y(n1955) );
  XOR2X1 U2302 ( .A(Inst_forkAE_KEY_INVERSE[106]), .B(
        Inst_forkAE_KEY_INVERSE[105]), .Y(n816) );
  XOR2X1 U2303 ( .A(n1794), .B(n1956), .Y(n1954) );
  XOR2X1 U2304 ( .A(n1059), .B(n1654), .Y(n1212) );
  XNOR2X1 U2305 ( .A(n1957), .B(n1958), .Y(n1059) );
  XOR2X1 U2306 ( .A(n179), .B(Inst_forkAE_KEY_INVERSE[155]), .Y(n1958) );
  XOR2X1 U2307 ( .A(n1959), .B(n1303), .Y(n1957) );
  XOR2X1 U2308 ( .A(Inst_forkAE_CURRENT_KEY_63_), .B(
        Inst_forkAE_KEY_INVERSE[90]), .Y(n1303) );
  OAI221X1 U2309 ( .A0(n1216), .A1(n1245), .B0(n1960), .B1(n1247), .C0(n1961), 
        .Y(Inst_forkAE_L_N16) );
  AOI22XL U2310 ( .A0(n1249), .A1(n1267), .B0(C1[14]), .B1(n135), .Y(n1961) );
  XOR2X1 U2311 ( .A(n1480), .B(n1962), .Y(n1267) );
  CLKINVX1 U2312 ( .A(n1675), .Y(n1962) );
  XNOR2X1 U2313 ( .A(n1963), .B(n1964), .Y(n1480) );
  XOR2X1 U2314 ( .A(n1965), .B(n1966), .Y(n1964) );
  XOR2X1 U2315 ( .A(Inst_forkAE_KEY_INVERSE[42]), .B(
        Inst_forkAE_KEY_INVERSE[170]), .Y(n1966) );
  XOR2X1 U2316 ( .A(n179), .B(Inst_forkAE_KEY_INVERSE[43]), .Y(n1965) );
  XOR2X1 U2317 ( .A(n1967), .B(n1968), .Y(n1963) );
  XOR2X1 U2318 ( .A(Inst_forkAE_KEY_INVERSE[105]), .B(n827), .Y(n1968) );
  XNOR2X1 U2319 ( .A(n1794), .B(n1969), .Y(n1967) );
  XOR2X1 U2320 ( .A(n131), .B(n1768), .Y(n1794) );
  CLKINVX1 U2321 ( .A(n1213), .Y(n1960) );
  XOR2X1 U2322 ( .A(n1064), .B(n1970), .Y(n1213) );
  CLKINVX1 U2323 ( .A(n1667), .Y(n1970) );
  XOR2X1 U2324 ( .A(n1971), .B(n1972), .Y(n1064) );
  XOR2X1 U2325 ( .A(Inst_forkAE_KEY_INVERSE[154]), .B(Inst_forkAE_CONST_ENC_2_), .Y(n1972) );
  XOR2X1 U2326 ( .A(n1973), .B(n1306), .Y(n1971) );
  XOR2X1 U2327 ( .A(Inst_forkAE_KEY_INVERSE[27]), .B(
        Inst_forkAE_KEY_INVERSE[89]), .Y(n1306) );
  OAI221X1 U2328 ( .A0(n1974), .A1(n1245), .B0(n1274), .B1(n1247), .C0(n1975), 
        .Y(Inst_forkAE_L_N15) );
  AOI22XL U2329 ( .A0(n1249), .A1(n1275), .B0(C1[13]), .B1(n135), .Y(n1975) );
  XOR2X1 U2330 ( .A(n1483), .B(n1976), .Y(n1275) );
  CLKINVX1 U2331 ( .A(n1687), .Y(n1976) );
  XOR2X1 U2332 ( .A(n1977), .B(C1[22]), .Y(n1687) );
  OR2X1 U2333 ( .A(C1[21]), .B(n1949), .Y(n1977) );
  CLKINVX1 U2334 ( .A(n1661), .Y(n1949) );
  XNOR2X1 U2335 ( .A(n1978), .B(n1979), .Y(n1483) );
  XOR2X1 U2336 ( .A(n1980), .B(n1981), .Y(n1979) );
  XOR2X1 U2337 ( .A(Inst_forkAE_CONST_ENC_2_), .B(C1[62]), .Y(n1981) );
  XOR2X1 U2338 ( .A(n181), .B(Inst_forkAE_KEY_INVERSE[169]), .Y(n1980) );
  XOR2X1 U2339 ( .A(n1982), .B(n827), .Y(n1978) );
  XOR2X1 U2340 ( .A(Inst_forkAE_KEY_INVERSE[104]), .B(
        Inst_forkAE_KEY_INVERSE[107]), .Y(n827) );
  XOR2X1 U2341 ( .A(n1983), .B(n454), .Y(n1982) );
  XOR2X1 U2342 ( .A(n578), .B(n573), .Y(n454) );
  CLKINVX1 U2343 ( .A(Inst_forkAE_KEY_INVERSE[42]), .Y(n573) );
  CLKINVX1 U2344 ( .A(Inst_forkAE_KEY_INVERSE[41]), .Y(n578) );
  CLKNAND2X2 U2345 ( .A(n1956), .B(n985), .Y(n1983) );
  CLKINVX1 U2346 ( .A(C1[61]), .Y(n985) );
  XNOR2X1 U2347 ( .A(n1067), .B(n1984), .Y(n1274) );
  CLKINVX1 U2348 ( .A(n1681), .Y(n1984) );
  XOR2X1 U2349 ( .A(n1985), .B(C0[22]), .Y(n1681) );
  NAND2BX1 U2350 ( .AN(C0[21]), .B(n1654), .Y(n1985) );
  XOR2X1 U2351 ( .A(n1986), .B(n1987), .Y(n1067) );
  XOR2X1 U2352 ( .A(C0[62]), .B(n1988), .Y(n1987) );
  XOR2X1 U2353 ( .A(Inst_forkAE_KEY_INVERSE[153]), .B(Inst_forkAE_CONST_ENC_1_), .Y(n1988) );
  XOR2X1 U2354 ( .A(n1989), .B(n1294), .Y(n1986) );
  XOR2X1 U2355 ( .A(Inst_forkAE_KEY_INVERSE[26]), .B(
        Inst_forkAE_KEY_INVERSE[88]), .Y(n1294) );
  NAND2BX1 U2356 ( .AN(C0[61]), .B(n1959), .Y(n1989) );
  OAI221X1 U2357 ( .A0(n1224), .A1(n1245), .B0(n1221), .B1(n1247), .C0(n1990), 
        .Y(Inst_forkAE_L_N14) );
  AOI22XL U2358 ( .A0(n1307), .A1(n1249), .B0(n135), .B1(C1[12]), .Y(n1990) );
  XOR2X1 U2359 ( .A(n1486), .B(n1991), .Y(n1307) );
  CLKINVX1 U2360 ( .A(n1706), .Y(n1991) );
  XOR2X1 U2361 ( .A(n1992), .B(C1[21]), .Y(n1706) );
  CLKNAND2X2 U2362 ( .A(n1675), .B(n1661), .Y(n1992) );
  XNOR2X1 U2363 ( .A(C1[20]), .B(n1993), .Y(n1661) );
  NOR2X1 U2364 ( .A(C1[22]), .B(C1[23]), .Y(n1993) );
  XOR2X1 U2365 ( .A(n1171), .B(n1994), .Y(n1675) );
  NOR2X1 U2366 ( .A(C1[21]), .B(C1[22]), .Y(n1994) );
  CLKINVX1 U2367 ( .A(C1[23]), .Y(n1171) );
  XOR2X1 U2368 ( .A(n1995), .B(n1996), .Y(n1486) );
  XOR2X1 U2369 ( .A(n1997), .B(n1998), .Y(n1996) );
  XOR2X1 U2370 ( .A(Inst_forkAE_KEY_INVERSE[168]), .B(
        Inst_forkAE_KEY_INVERSE[107]), .Y(n1998) );
  XOR2X1 U2371 ( .A(Inst_forkAE_KEY_INVERSE[41]), .B(
        Inst_forkAE_KEY_INVERSE[40]), .Y(n1997) );
  XOR2X1 U2372 ( .A(n1999), .B(n2000), .Y(n1995) );
  XOR2X1 U2373 ( .A(n2001), .B(C1[61]), .Y(n1999) );
  NAND2BX1 U2374 ( .AN(n1969), .B(n1956), .Y(n2001) );
  XNOR2X1 U2375 ( .A(C1[60]), .B(n2002), .Y(n1956) );
  NOR2X1 U2376 ( .A(C1[62]), .B(C1[63]), .Y(n2002) );
  XNOR2X1 U2377 ( .A(n976), .B(n2003), .Y(n1969) );
  NOR2X1 U2378 ( .A(C1[61]), .B(C1[62]), .Y(n2003) );
  CLKINVX1 U2379 ( .A(C1[63]), .Y(n976) );
  XOR2X1 U2380 ( .A(n1071), .B(n1696), .Y(n1221) );
  XNOR2X1 U2381 ( .A(n2004), .B(C0[21]), .Y(n1696) );
  CLKNAND2X2 U2382 ( .A(n1667), .B(n1654), .Y(n2004) );
  XNOR2X1 U2383 ( .A(C0[20]), .B(n2005), .Y(n1654) );
  NOR2X1 U2384 ( .A(C0[22]), .B(C0[23]), .Y(n2005) );
  XNOR2X1 U2385 ( .A(C0[23]), .B(n2006), .Y(n1667) );
  NOR2X1 U2386 ( .A(C0[21]), .B(C0[22]), .Y(n2006) );
  XOR2X1 U2387 ( .A(n2007), .B(n2008), .Y(n1071) );
  XNOR2X1 U2388 ( .A(n1299), .B(n1768), .Y(n2008) );
  XOR2X1 U2389 ( .A(Inst_forkAE_CURRENT_KEY_124_), .B(
        Inst_forkAE_KEY_INVERSE[25]), .Y(n1299) );
  XOR2X1 U2390 ( .A(n2009), .B(n2010), .Y(n2007) );
  XOR2X1 U2391 ( .A(Inst_forkAE_KEY_INVERSE[152]), .B(C0[61]), .Y(n2010) );
  CLKNAND2X2 U2392 ( .A(n1973), .B(n1959), .Y(n2009) );
  XNOR2X1 U2393 ( .A(C0[60]), .B(n2011), .Y(n1959) );
  NOR2X1 U2394 ( .A(C0[62]), .B(C0[63]), .Y(n2011) );
  XNOR2X1 U2395 ( .A(C0[63]), .B(n2012), .Y(n1973) );
  NOR2X1 U2396 ( .A(C0[61]), .B(C0[62]), .Y(n2012) );
  XOR2X1 U2397 ( .A(n2013), .B(n2014), .Y(n1224) );
  CLKNAND2X2 U2398 ( .A(n1211), .B(n1216), .Y(n2013) );
  XOR2X1 U2399 ( .A(n2015), .B(n2016), .Y(n1211) );
  CLKNAND2X2 U2400 ( .A(n1216), .B(n1974), .Y(n2015) );
  XOR2X1 U2401 ( .A(n2017), .B(n2018), .Y(n1216) );
  XOR2X1 U2402 ( .A(C0[49]), .B(C0[1]), .Y(n2018) );
  OR2X1 U2403 ( .A(n2014), .B(n1219), .Y(n2017) );
  CLKINVX1 U2404 ( .A(n1974), .Y(n1219) );
  XOR2X1 U2405 ( .A(n2019), .B(n2020), .Y(n1974) );
  NOR2X1 U2406 ( .A(n2014), .B(n2016), .Y(n2020) );
  XOR2X1 U2407 ( .A(C0[2]), .B(C0[50]), .Y(n2016) );
  XNOR2X1 U2408 ( .A(C0[0]), .B(C0[48]), .Y(n2019) );
  XOR2X1 U2409 ( .A(C0[51]), .B(C0[3]), .Y(n2014) );
  OAI221X1 U2410 ( .A0(n1228), .A1(n1245), .B0(n2021), .B1(n1247), .C0(n2022), 
        .Y(Inst_forkAE_L_N13) );
  AOI22XL U2411 ( .A0(n1249), .A1(n1315), .B0(C1[11]), .B1(n135), .Y(n2022) );
  XOR2X1 U2412 ( .A(n1515), .B(n2023), .Y(n1315) );
  XNOR2X1 U2413 ( .A(n2024), .B(n2025), .Y(n1515) );
  XOR2X1 U2414 ( .A(Inst_forkAE_KEY_INVERSE[102]), .B(n2026), .Y(n2025) );
  XOR2X1 U2415 ( .A(Inst_forkAE_KEY_INVERSE[36]), .B(
        Inst_forkAE_KEY_INVERSE[167]), .Y(n2026) );
  XNOR2X1 U2416 ( .A(n2027), .B(n2028), .Y(n2024) );
  CLKINVX1 U2417 ( .A(n1225), .Y(n2021) );
  XNOR2X1 U2418 ( .A(n1076), .B(n1727), .Y(n1225) );
  XNOR2X1 U2419 ( .A(n2029), .B(n2030), .Y(n1076) );
  XNOR2X1 U2420 ( .A(Inst_forkAE_KEY_INVERSE[131]), .B(n1360), .Y(n2029) );
  XOR2X1 U2421 ( .A(Inst_forkAE_CURRENT_KEY_59_), .B(
        Inst_forkAE_KEY_INVERSE[66]), .Y(n1360) );
  OAI221X1 U2422 ( .A0(n1232), .A1(n1245), .B0(n1320), .B1(n1247), .C0(n2031), 
        .Y(Inst_forkAE_L_N12) );
  AOI22XL U2423 ( .A0(n1249), .A1(n1321), .B0(C1[10]), .B1(n135), .Y(n2031) );
  XNOR2X1 U2424 ( .A(n1518), .B(n1745), .Y(n1321) );
  XNOR2X1 U2425 ( .A(n2032), .B(n2033), .Y(n1518) );
  XOR2X1 U2426 ( .A(Inst_forkAE_KEY_INVERSE[166]), .B(n2034), .Y(n2033) );
  XOR2X1 U2427 ( .A(Inst_forkAE_KEY_INVERSE[39]), .B(
        Inst_forkAE_KEY_INVERSE[38]), .Y(n2034) );
  XNOR2X1 U2428 ( .A(n2027), .B(n2035), .Y(n2032) );
  XOR2X1 U2429 ( .A(n602), .B(n854), .Y(n2027) );
  CLKINVX1 U2430 ( .A(Inst_forkAE_KEY_INVERSE[101]), .Y(n602) );
  XOR2X1 U2431 ( .A(n1080), .B(n1739), .Y(n1320) );
  XNOR2X1 U2432 ( .A(n2036), .B(n2037), .Y(n1080) );
  XNOR2X1 U2433 ( .A(Inst_forkAE_KEY_INVERSE[130]), .B(n1362), .Y(n2036) );
  XOR2X1 U2434 ( .A(Inst_forkAE_KEY_INVERSE[3]), .B(
        Inst_forkAE_KEY_INVERSE[65]), .Y(n1362) );
  OAI221X1 U2435 ( .A0(n2038), .A1(n1245), .B0(n1234), .B1(n1247), .C0(n2039), 
        .Y(Inst_forkAE_L_N11) );
  AOI22XL U2436 ( .A0(n1249), .A1(n1338), .B0(n135), .B1(C1[9]), .Y(n2039) );
  XOR2X1 U2437 ( .A(n1521), .B(n2040), .Y(n1338) );
  CLKINVX1 U2438 ( .A(n1769), .Y(n2040) );
  XOR2X1 U2439 ( .A(n2041), .B(C1[18]), .Y(n1769) );
  OR2X1 U2440 ( .A(C1[17]), .B(n2023), .Y(n2041) );
  CLKINVX1 U2441 ( .A(n1734), .Y(n2023) );
  XNOR2X1 U2442 ( .A(n2042), .B(n2043), .Y(n1521) );
  XOR2X1 U2443 ( .A(n485), .B(n854), .Y(n2043) );
  XOR2X1 U2444 ( .A(Inst_forkAE_KEY_INVERSE[100]), .B(
        Inst_forkAE_KEY_INVERSE[103]), .Y(n854) );
  XNOR2X1 U2445 ( .A(n204), .B(Inst_forkAE_KEY_INVERSE[38]), .Y(n485) );
  CLKINVX1 U2446 ( .A(Inst_forkAE_KEY_INVERSE[37]), .Y(n204) );
  XOR2X1 U2447 ( .A(n2044), .B(n2045), .Y(n2042) );
  XOR2X1 U2448 ( .A(Inst_forkAE_KEY_INVERSE[165]), .B(C1[58]), .Y(n2045) );
  NAND2BX1 U2449 ( .AN(C1[57]), .B(n2028), .Y(n2044) );
  XOR2X1 U2450 ( .A(n1084), .B(n1758), .Y(n1234) );
  XNOR2X1 U2451 ( .A(n2046), .B(C0[18]), .Y(n1758) );
  NAND2BX1 U2452 ( .AN(C0[17]), .B(n1727), .Y(n2046) );
  XOR2X1 U2453 ( .A(n2047), .B(n2048), .Y(n1084) );
  XOR2X1 U2454 ( .A(Inst_forkAE_KEY_INVERSE[129]), .B(C0[58]), .Y(n2048) );
  XOR2X1 U2455 ( .A(n2049), .B(n1354), .Y(n2047) );
  XOR2X1 U2456 ( .A(Inst_forkAE_KEY_INVERSE[2]), .B(
        Inst_forkAE_KEY_INVERSE[64]), .Y(n1354) );
  NAND2BX1 U2457 ( .AN(C0[57]), .B(n2030), .Y(n2049) );
  OAI221X1 U2458 ( .A0(n1241), .A1(n1245), .B0(n1238), .B1(n1247), .C0(n2050), 
        .Y(Inst_forkAE_L_N10) );
  AOI22XL U2459 ( .A0(n1249), .A1(n1363), .B0(n135), .B1(C1[8]), .Y(n2050) );
  XOR2X1 U2460 ( .A(n1523), .B(n2051), .Y(n1363) );
  CLKINVX1 U2461 ( .A(n1797), .Y(n2051) );
  XOR2X1 U2462 ( .A(n2052), .B(C1[17]), .Y(n1797) );
  CLKNAND2X2 U2463 ( .A(n1745), .B(n1734), .Y(n2052) );
  XNOR2X1 U2464 ( .A(C1[16]), .B(n2053), .Y(n1734) );
  NOR2X1 U2465 ( .A(C1[18]), .B(C1[19]), .Y(n2053) );
  XNOR2X1 U2466 ( .A(C1[19]), .B(n2054), .Y(n1745) );
  NOR2X1 U2467 ( .A(C1[17]), .B(C1[18]), .Y(n2054) );
  XNOR2X1 U2468 ( .A(n2055), .B(n2056), .Y(n1523) );
  XOR2X1 U2469 ( .A(Inst_forkAE_KEY_INVERSE[164]), .B(n2057), .Y(n2056) );
  XOR2X1 U2470 ( .A(Inst_forkAE_KEY_INVERSE[37]), .B(
        Inst_forkAE_KEY_INVERSE[36]), .Y(n2057) );
  XOR2X1 U2471 ( .A(n2058), .B(n2059), .Y(n2055) );
  XOR2X1 U2472 ( .A(Inst_forkAE_KEY_INVERSE[103]), .B(C1[57]), .Y(n2059) );
  CLKNAND2X2 U2473 ( .A(n2035), .B(n2028), .Y(n2058) );
  XNOR2X1 U2474 ( .A(C1[56]), .B(n2060), .Y(n2028) );
  NOR2X1 U2475 ( .A(C1[58]), .B(C1[59]), .Y(n2060) );
  XNOR2X1 U2476 ( .A(C1[59]), .B(n2061), .Y(n2035) );
  NOR2X1 U2477 ( .A(C1[57]), .B(C1[58]), .Y(n2061) );
  CLKNAND2X2 U2478 ( .A(n184), .B(n1257), .Y(n1247) );
  AOI31X1 U2479 ( .A0(n2062), .A1(n180), .A2(n2063), .B0(n2064), .Y(n1249) );
  NOR3X1 U2480 ( .A(n185), .B(n183), .C(n2065), .Y(n2062) );
  CLKINVX1 U2481 ( .A(Inst_forkAE_CONST_ENC_5_), .Y(n183) );
  XOR2X1 U2482 ( .A(n1089), .B(n2066), .Y(n1238) );
  CLKINVX1 U2483 ( .A(n1777), .Y(n2066) );
  XOR2X1 U2484 ( .A(n2067), .B(C0[17]), .Y(n1777) );
  CLKNAND2X2 U2485 ( .A(n1739), .B(n1727), .Y(n2067) );
  XNOR2X1 U2486 ( .A(C0[16]), .B(n2068), .Y(n1727) );
  NOR2X1 U2487 ( .A(C0[18]), .B(C0[19]), .Y(n2068) );
  XNOR2X1 U2488 ( .A(C0[19]), .B(n2069), .Y(n1739) );
  NOR2X1 U2489 ( .A(C0[17]), .B(C0[18]), .Y(n2069) );
  XOR2X1 U2490 ( .A(n2070), .B(n2071), .Y(n1089) );
  XOR2X1 U2491 ( .A(Inst_forkAE_KEY_INVERSE[128]), .B(C0[57]), .Y(n2071) );
  XOR2X1 U2492 ( .A(n2072), .B(n1358), .Y(n2070) );
  XOR2X1 U2493 ( .A(Inst_forkAE_CURRENT_KEY_120_), .B(
        Inst_forkAE_KEY_INVERSE[1]), .Y(n1358) );
  CLKNAND2X2 U2494 ( .A(n2037), .B(n2030), .Y(n2072) );
  XNOR2X1 U2495 ( .A(C0[56]), .B(n2073), .Y(n2030) );
  NOR2X1 U2496 ( .A(C0[58]), .B(C0[59]), .Y(n2073) );
  XNOR2X1 U2497 ( .A(C0[59]), .B(n2074), .Y(n2037) );
  NOR2X1 U2498 ( .A(C0[57]), .B(C0[58]), .Y(n2074) );
  NOR3BX1 U2499 ( .AN(n2075), .B(n184), .C(n1243), .Y(n1251) );
  NAND4X1 U2500 ( .A(Inst_forkAE_CONST_ENC_1_), .B(Inst_forkAE_CONST_ENC_2_), 
        .C(n181), .D(n2076), .Y(n2075) );
  NOR4X1 U2501 ( .A(n180), .B(n179), .C(Inst_forkAE_CONST_ENC_5_), .D(n182), 
        .Y(n2076) );
  CLKINVX1 U2502 ( .A(Inst_forkAE_CONST_DEC_6_), .Y(n182) );
  XOR2X1 U2503 ( .A(n2077), .B(n2078), .Y(n1241) );
  CLKNAND2X2 U2504 ( .A(n1228), .B(n1232), .Y(n2077) );
  XOR2X1 U2505 ( .A(n2079), .B(n2080), .Y(n1228) );
  CLKNAND2X2 U2506 ( .A(n1232), .B(n2038), .Y(n2079) );
  XOR2X1 U2507 ( .A(n2081), .B(n2082), .Y(n1232) );
  XOR2X1 U2508 ( .A(C0[61]), .B(C0[13]), .Y(n2082) );
  OR2X1 U2509 ( .A(n2078), .B(n1236), .Y(n2081) );
  CLKINVX1 U2510 ( .A(n2038), .Y(n1236) );
  XOR2X1 U2511 ( .A(n2083), .B(n2084), .Y(n2038) );
  NOR2X1 U2512 ( .A(n2078), .B(n2080), .Y(n2084) );
  XOR2X1 U2513 ( .A(C0[14]), .B(C0[62]), .Y(n2080) );
  XNOR2X1 U2514 ( .A(C0[12]), .B(C0[60]), .Y(n2083) );
  XOR2X1 U2515 ( .A(C0[63]), .B(C0[15]), .Y(n2078) );
  CLKNAND2X2 U2516 ( .A(n2085), .B(n951), .Y(Inst_forkAE_FSM_X_N43) );
  CLKNAND2X2 U2517 ( .A(Inst_forkAE_FSM_X_state_1_), .B(n957), .Y(n951) );
  MXI2X1 U2518 ( .A(n2086), .B(n2087), .S0(n2088), .Y(n2085) );
  NOR3X1 U2519 ( .A(n957), .B(Inst_forkAE_FSM_X_state_1_), .C(n958), .Y(n2086)
         );
  CLKINVX1 U2520 ( .A(Inst_forkAE_FSM_X_state_2_), .Y(n958) );
  OAI2B2X1 U2521 ( .A1N(n2087), .A0(n957), .B0(n2089), .B1(n1244), .Y(
        Inst_forkAE_FSM_X_N42) );
  AOI21X1 U2522 ( .A0(GO), .A1(ENC_DEC_MODE), .B0(Inst_forkAE_FSM_X_state_2_), 
        .Y(n2089) );
  OAI31X1 U2523 ( .A0(n950), .A1(ENC_DEC_MODE), .A2(n1244), .B0(n2090), .Y(
        Inst_forkAE_FSM_X_N41) );
  MXI2X1 U2524 ( .A(Inst_forkAE_FSM_X_state_2_), .B(n2091), .S0(
        Inst_forkAE_FSM_X_state_0_), .Y(n2090) );
  AOI21X1 U2525 ( .A0(Inst_forkAE_FSM_X_state_1_), .A1(
        Inst_forkAE_FSM_X_state_2_), .B0(n2088), .Y(n2091) );
  MXI2X1 U2526 ( .A(n2092), .B(n2093), .S0(n2064), .Y(n2088) );
  NAND2BX1 U2527 ( .AN(n2094), .B(Inst_forkAE_CONST_ENC_2_), .Y(n2093) );
  CLKNAND2X2 U2528 ( .A(n957), .B(n956), .Y(n1244) );
  CLKINVX1 U2529 ( .A(GO), .Y(n950) );
  NOR2X1 U2530 ( .A(n2095), .B(n2096), .Y(Inst_forkAE_ConstGen_N30) );
  MXI2X1 U2531 ( .A(n2097), .B(n131), .S0(n184), .Y(n2096) );
  CLKNAND2X2 U2532 ( .A(Inst_forkAE_FSM_X_state_0_), .B(n2098), .Y(n2097) );
  XOR2X1 U2533 ( .A(Inst_forkAE_CONST_ENC_1_), .B(Inst_forkAE_CONST_DEC_6_), 
        .Y(n2098) );
  AOI21X1 U2534 ( .A0(n2099), .A1(n2100), .B0(n2095), .Y(
        Inst_forkAE_ConstGen_N28) );
  MXI2X1 U2535 ( .A(n131), .B(n133), .S0(n184), .Y(n2099) );
  AOI21X1 U2536 ( .A0(n2101), .A1(n2100), .B0(n2095), .Y(
        Inst_forkAE_ConstGen_N25) );
  NOR2X1 U2537 ( .A(n2064), .B(Inst_forkAE_FSM_X_state_0_), .Y(n2095) );
  MXI2X1 U2538 ( .A(n132), .B(Inst_forkAE_CONST_ENC_1_), .S0(n184), .Y(n2101)
         );
  CLKNAND2X2 U2539 ( .A(n2102), .B(n2100), .Y(Inst_forkAE_ConstGen_N24) );
  CLKNAND2X2 U2540 ( .A(n2064), .B(n957), .Y(n2100) );
  MXI2X1 U2541 ( .A(Inst_forkAE_CONST_ENC_2_), .B(n2103), .S0(n184), .Y(n2102)
         );
  NOR2X1 U2542 ( .A(n1768), .B(n957), .Y(n2103) );
  MX2X1 U2543 ( .A(IDtReg[48]), .B(IDt[48]), .S0(ld_rec), .Y(Inst_RegIDt_n99)
         );
  MX2X1 U2544 ( .A(IDtReg[47]), .B(IDt[47]), .S0(ld_rec), .Y(Inst_RegIDt_n97)
         );
  MX2X1 U2545 ( .A(IDtReg[46]), .B(IDt[46]), .S0(ld_rec), .Y(Inst_RegIDt_n95)
         );
  MX2X1 U2546 ( .A(IDtReg[45]), .B(IDt[45]), .S0(ld_rec), .Y(Inst_RegIDt_n93)
         );
  MX2X1 U2547 ( .A(IDtReg[44]), .B(IDt[44]), .S0(ld_rec), .Y(Inst_RegIDt_n91)
         );
  MX2X1 U2548 ( .A(IDtReg[3]), .B(IDt[3]), .S0(ld_rec), .Y(Inst_RegIDt_n9) );
  MX2X1 U2549 ( .A(IDtReg[43]), .B(IDt[43]), .S0(ld_rec), .Y(Inst_RegIDt_n89)
         );
  MX2X1 U2550 ( .A(IDtReg[42]), .B(IDt[42]), .S0(ld_rec), .Y(Inst_RegIDt_n87)
         );
  MX2X1 U2551 ( .A(IDtReg[41]), .B(IDt[41]), .S0(ld_rec), .Y(Inst_RegIDt_n85)
         );
  MX2X1 U2552 ( .A(IDtReg[40]), .B(IDt[40]), .S0(ld_rec), .Y(Inst_RegIDt_n83)
         );
  MX2X1 U2553 ( .A(IDtReg[39]), .B(IDt[39]), .S0(ld_rec), .Y(Inst_RegIDt_n81)
         );
  MX2X1 U2554 ( .A(IDtReg[38]), .B(IDt[38]), .S0(ld_rec), .Y(Inst_RegIDt_n79)
         );
  MX2X1 U2555 ( .A(IDtReg[37]), .B(IDt[37]), .S0(ld_rec), .Y(Inst_RegIDt_n77)
         );
  MX2X1 U2556 ( .A(IDtReg[36]), .B(IDt[36]), .S0(ld_rec), .Y(Inst_RegIDt_n75)
         );
  MX2X1 U2557 ( .A(IDtReg[35]), .B(IDt[35]), .S0(ld_rec), .Y(Inst_RegIDt_n73)
         );
  MX2X1 U2558 ( .A(IDtReg[34]), .B(IDt[34]), .S0(ld_rec), .Y(Inst_RegIDt_n71)
         );
  MX2X1 U2559 ( .A(IDtReg[2]), .B(IDt[2]), .S0(ld_rec), .Y(Inst_RegIDt_n7) );
  MX2X1 U2560 ( .A(IDtReg[33]), .B(IDt[33]), .S0(ld_rec), .Y(Inst_RegIDt_n69)
         );
  MX2X1 U2561 ( .A(IDtReg[32]), .B(IDt[32]), .S0(ld_rec), .Y(Inst_RegIDt_n67)
         );
  MX2X1 U2562 ( .A(IDtReg[31]), .B(IDt[31]), .S0(ld_rec), .Y(Inst_RegIDt_n65)
         );
  MX2X1 U2563 ( .A(IDtReg[30]), .B(IDt[30]), .S0(ld_rec), .Y(Inst_RegIDt_n63)
         );
  MX2X1 U2564 ( .A(IDtReg[29]), .B(IDt[29]), .S0(ld_rec), .Y(Inst_RegIDt_n61)
         );
  MX2X1 U2565 ( .A(IDtReg[28]), .B(IDt[28]), .S0(ld_rec), .Y(Inst_RegIDt_n59)
         );
  MX2X1 U2566 ( .A(IDtReg[27]), .B(IDt[27]), .S0(ld_rec), .Y(Inst_RegIDt_n57)
         );
  MX2X1 U2567 ( .A(IDtReg[26]), .B(IDt[26]), .S0(ld_rec), .Y(Inst_RegIDt_n55)
         );
  MX2X1 U2568 ( .A(IDtReg[25]), .B(IDt[25]), .S0(ld_rec), .Y(Inst_RegIDt_n53)
         );
  MX2X1 U2569 ( .A(IDtReg[24]), .B(IDt[24]), .S0(ld_rec), .Y(Inst_RegIDt_n51)
         );
  MX2X1 U2570 ( .A(IDtReg[1]), .B(IDt[1]), .S0(ld_rec), .Y(Inst_RegIDt_n5) );
  MX2X1 U2571 ( .A(IDtReg[23]), .B(IDt[23]), .S0(ld_rec), .Y(Inst_RegIDt_n49)
         );
  MX2X1 U2572 ( .A(IDtReg[22]), .B(IDt[22]), .S0(ld_rec), .Y(Inst_RegIDt_n47)
         );
  MX2X1 U2573 ( .A(IDtReg[21]), .B(IDt[21]), .S0(ld_rec), .Y(Inst_RegIDt_n45)
         );
  MX2X1 U2574 ( .A(IDtReg[20]), .B(IDt[20]), .S0(ld_rec), .Y(Inst_RegIDt_n43)
         );
  MX2X1 U2575 ( .A(IDtReg[19]), .B(IDt[19]), .S0(ld_rec), .Y(Inst_RegIDt_n41)
         );
  MX2X1 U2576 ( .A(IDtReg[18]), .B(IDt[18]), .S0(ld_rec), .Y(Inst_RegIDt_n39)
         );
  MX2X1 U2577 ( .A(IDtReg[17]), .B(IDt[17]), .S0(ld_rec), .Y(Inst_RegIDt_n37)
         );
  MX2X1 U2578 ( .A(IDtReg[16]), .B(IDt[16]), .S0(ld_rec), .Y(Inst_RegIDt_n35)
         );
  MX2X1 U2579 ( .A(IDtReg[15]), .B(IDt[15]), .S0(ld_rec), .Y(Inst_RegIDt_n33)
         );
  MX2X1 U2580 ( .A(IDtReg[14]), .B(IDt[14]), .S0(ld_rec), .Y(Inst_RegIDt_n31)
         );
  MX2X1 U2581 ( .A(IDtReg[0]), .B(IDt[0]), .S0(ld_rec), .Y(Inst_RegIDt_n3) );
  MX2X1 U2582 ( .A(IDtReg[13]), .B(IDt[13]), .S0(ld_rec), .Y(Inst_RegIDt_n29)
         );
  MX2X1 U2583 ( .A(IDtReg[12]), .B(IDt[12]), .S0(ld_rec), .Y(Inst_RegIDt_n27)
         );
  MX2X1 U2584 ( .A(IDtReg[11]), .B(IDt[11]), .S0(ld_rec), .Y(Inst_RegIDt_n25)
         );
  MX2X1 U2585 ( .A(IDtReg[10]), .B(IDt[10]), .S0(ld_rec), .Y(Inst_RegIDt_n23)
         );
  MX2X1 U2586 ( .A(IDtReg[9]), .B(IDt[9]), .S0(ld_rec), .Y(Inst_RegIDt_n21) );
  MX2X1 U2587 ( .A(IDtReg[8]), .B(IDt[8]), .S0(ld_rec), .Y(Inst_RegIDt_n19) );
  MX2X1 U2588 ( .A(IDtReg[7]), .B(IDt[7]), .S0(ld_rec), .Y(Inst_RegIDt_n17) );
  MX2X1 U2589 ( .A(IDtReg[6]), .B(IDt[6]), .S0(ld_rec), .Y(Inst_RegIDt_n15) );
  MX2X1 U2590 ( .A(IDtReg[63]), .B(IDt[63]), .S0(ld_rec), .Y(Inst_RegIDt_n130)
         );
  MX2X1 U2591 ( .A(IDtReg[5]), .B(IDt[5]), .S0(ld_rec), .Y(Inst_RegIDt_n13) );
  MX2X1 U2592 ( .A(IDtReg[62]), .B(IDt[62]), .S0(ld_rec), .Y(Inst_RegIDt_n127)
         );
  MX2X1 U2593 ( .A(IDtReg[61]), .B(IDt[61]), .S0(ld_rec), .Y(Inst_RegIDt_n125)
         );
  MX2X1 U2594 ( .A(IDtReg[60]), .B(IDt[60]), .S0(ld_rec), .Y(Inst_RegIDt_n123)
         );
  MX2X1 U2595 ( .A(IDtReg[59]), .B(IDt[59]), .S0(ld_rec), .Y(Inst_RegIDt_n121)
         );
  MX2X1 U2596 ( .A(IDtReg[58]), .B(IDt[58]), .S0(ld_rec), .Y(Inst_RegIDt_n119)
         );
  MX2X1 U2597 ( .A(IDtReg[57]), .B(IDt[57]), .S0(ld_rec), .Y(Inst_RegIDt_n117)
         );
  MX2X1 U2598 ( .A(IDtReg[56]), .B(IDt[56]), .S0(ld_rec), .Y(Inst_RegIDt_n115)
         );
  MX2X1 U2599 ( .A(IDtReg[55]), .B(IDt[55]), .S0(ld_rec), .Y(Inst_RegIDt_n113)
         );
  MX2X1 U2600 ( .A(IDtReg[54]), .B(IDt[54]), .S0(ld_rec), .Y(Inst_RegIDt_n111)
         );
  MX2X1 U2601 ( .A(IDtReg[4]), .B(IDt[4]), .S0(ld_rec), .Y(Inst_RegIDt_n11) );
  MX2X1 U2602 ( .A(IDtReg[53]), .B(IDt[53]), .S0(ld_rec), .Y(Inst_RegIDt_n109)
         );
  MX2X1 U2603 ( .A(IDtReg[52]), .B(IDt[52]), .S0(ld_rec), .Y(Inst_RegIDt_n107)
         );
  MX2X1 U2604 ( .A(IDtReg[51]), .B(IDt[51]), .S0(ld_rec), .Y(Inst_RegIDt_n105)
         );
  MX2X1 U2605 ( .A(IDtReg[50]), .B(IDt[50]), .S0(ld_rec), .Y(Inst_RegIDt_n103)
         );
  MX2X1 U2606 ( .A(IDtReg[49]), .B(IDt[49]), .S0(ld_rec), .Y(Inst_RegIDt_n101)
         );
  MX2X1 U2607 ( .A(IDstReg[48]), .B(IDst[48]), .S0(ld_rec), .Y(n2718) );
  MX2X1 U2608 ( .A(IDstReg[47]), .B(IDst[47]), .S0(ld_rec), .Y(n2716) );
  MX2X1 U2609 ( .A(IDstReg[46]), .B(IDst[46]), .S0(ld_rec), .Y(n2714) );
  MX2X1 U2610 ( .A(IDstReg[45]), .B(IDst[45]), .S0(ld_rec), .Y(n2712) );
  MX2X1 U2611 ( .A(IDstReg[44]), .B(IDst[44]), .S0(ld_rec), .Y(n2710) );
  MX2X1 U2612 ( .A(IDstReg[3]), .B(IDst[3]), .S0(ld_rec), .Y(n2628) );
  MX2X1 U2613 ( .A(IDstReg[43]), .B(IDst[43]), .S0(ld_rec), .Y(n2708) );
  MX2X1 U2614 ( .A(IDstReg[42]), .B(IDst[42]), .S0(ld_rec), .Y(n2706) );
  MX2X1 U2615 ( .A(IDstReg[41]), .B(IDst[41]), .S0(ld_rec), .Y(n2704) );
  MX2X1 U2616 ( .A(IDstReg[40]), .B(IDst[40]), .S0(ld_rec), .Y(n2702) );
  MX2X1 U2617 ( .A(IDstReg[39]), .B(IDst[39]), .S0(ld_rec), .Y(n2700) );
  MX2X1 U2618 ( .A(IDstReg[38]), .B(IDst[38]), .S0(ld_rec), .Y(n2698) );
  MX2X1 U2619 ( .A(IDstReg[37]), .B(IDst[37]), .S0(ld_rec), .Y(n2696) );
  MX2X1 U2620 ( .A(IDstReg[36]), .B(IDst[36]), .S0(ld_rec), .Y(n2694) );
  MX2X1 U2621 ( .A(IDstReg[35]), .B(IDst[35]), .S0(ld_rec), .Y(n2692) );
  MX2X1 U2622 ( .A(IDstReg[34]), .B(IDst[34]), .S0(ld_rec), .Y(n2690) );
  MX2X1 U2623 ( .A(IDstReg[2]), .B(IDst[2]), .S0(ld_rec), .Y(n2626) );
  MX2X1 U2624 ( .A(IDstReg[33]), .B(IDst[33]), .S0(ld_rec), .Y(n2688) );
  MX2X1 U2625 ( .A(IDstReg[32]), .B(IDst[32]), .S0(ld_rec), .Y(n2686) );
  MX2X1 U2626 ( .A(IDstReg[31]), .B(IDst[31]), .S0(ld_rec), .Y(n2684) );
  MX2X1 U2627 ( .A(IDstReg[30]), .B(IDst[30]), .S0(ld_rec), .Y(n2682) );
  MX2X1 U2628 ( .A(IDstReg[29]), .B(IDst[29]), .S0(ld_rec), .Y(n2680) );
  MX2X1 U2629 ( .A(IDstReg[28]), .B(IDst[28]), .S0(ld_rec), .Y(n2678) );
  MX2X1 U2630 ( .A(IDstReg[27]), .B(IDst[27]), .S0(ld_rec), .Y(n2676) );
  MX2X1 U2631 ( .A(IDstReg[26]), .B(IDst[26]), .S0(ld_rec), .Y(n2674) );
  MX2X1 U2632 ( .A(IDstReg[25]), .B(IDst[25]), .S0(ld_rec), .Y(n2672) );
  MX2X1 U2633 ( .A(IDstReg[24]), .B(IDst[24]), .S0(ld_rec), .Y(n2670) );
  MX2X1 U2634 ( .A(IDstReg[1]), .B(IDst[1]), .S0(ld_rec), .Y(n2624) );
  MX2X1 U2635 ( .A(IDstReg[23]), .B(IDst[23]), .S0(ld_rec), .Y(n2668) );
  MX2X1 U2636 ( .A(IDstReg[22]), .B(IDst[22]), .S0(ld_rec), .Y(n2666) );
  MX2X1 U2637 ( .A(IDstReg[21]), .B(IDst[21]), .S0(ld_rec), .Y(n2664) );
  MX2X1 U2638 ( .A(IDstReg[20]), .B(IDst[20]), .S0(ld_rec), .Y(n2662) );
  MX2X1 U2639 ( .A(IDstReg[19]), .B(IDst[19]), .S0(ld_rec), .Y(n2660) );
  MX2X1 U2640 ( .A(IDstReg[18]), .B(IDst[18]), .S0(ld_rec), .Y(n2658) );
  MX2X1 U2641 ( .A(IDstReg[17]), .B(IDst[17]), .S0(ld_rec), .Y(n2656) );
  MX2X1 U2642 ( .A(IDstReg[16]), .B(IDst[16]), .S0(ld_rec), .Y(n2654) );
  MX2X1 U2643 ( .A(IDstReg[15]), .B(IDst[15]), .S0(ld_rec), .Y(n2652) );
  MX2X1 U2644 ( .A(IDstReg[14]), .B(IDst[14]), .S0(ld_rec), .Y(n2650) );
  MX2X1 U2645 ( .A(IDstReg[0]), .B(IDst[0]), .S0(ld_rec), .Y(n2622) );
  MX2X1 U2646 ( .A(IDstReg[13]), .B(IDst[13]), .S0(ld_rec), .Y(n2648) );
  MX2X1 U2647 ( .A(IDstReg[12]), .B(IDst[12]), .S0(ld_rec), .Y(n2646) );
  MX2X1 U2648 ( .A(IDstReg[11]), .B(IDst[11]), .S0(ld_rec), .Y(n2644) );
  MX2X1 U2649 ( .A(IDstReg[10]), .B(IDst[10]), .S0(ld_rec), .Y(n2642) );
  MX2X1 U2650 ( .A(IDstReg[9]), .B(IDst[9]), .S0(ld_rec), .Y(n2640) );
  MX2X1 U2651 ( .A(IDstReg[8]), .B(IDst[8]), .S0(ld_rec), .Y(n2638) );
  MX2X1 U2652 ( .A(IDstReg[7]), .B(IDst[7]), .S0(ld_rec), .Y(n2636) );
  MX2X1 U2653 ( .A(IDstReg[6]), .B(IDst[6]), .S0(ld_rec), .Y(n2634) );
  MX2X1 U2654 ( .A(IDstReg[63]), .B(IDst[63]), .S0(ld_rec), .Y(n2748) );
  MX2X1 U2655 ( .A(IDstReg[5]), .B(IDst[5]), .S0(ld_rec), .Y(n2632) );
  MX2X1 U2656 ( .A(IDstReg[62]), .B(IDst[62]), .S0(ld_rec), .Y(n2746) );
  MX2X1 U2657 ( .A(IDstReg[61]), .B(IDst[61]), .S0(ld_rec), .Y(n2744) );
  MX2X1 U2658 ( .A(IDstReg[60]), .B(IDst[60]), .S0(ld_rec), .Y(n2742) );
  MX2X1 U2659 ( .A(IDstReg[59]), .B(IDst[59]), .S0(ld_rec), .Y(n2740) );
  MX2X1 U2660 ( .A(IDstReg[58]), .B(IDst[58]), .S0(ld_rec), .Y(n2738) );
  MX2X1 U2661 ( .A(IDstReg[57]), .B(IDst[57]), .S0(ld_rec), .Y(n2736) );
  MX2X1 U2662 ( .A(IDstReg[56]), .B(IDst[56]), .S0(ld_rec), .Y(n2734) );
  MX2X1 U2663 ( .A(IDstReg[55]), .B(IDst[55]), .S0(ld_rec), .Y(n2732) );
  MX2X1 U2664 ( .A(IDstReg[54]), .B(IDst[54]), .S0(ld_rec), .Y(n2730) );
  MX2X1 U2665 ( .A(IDstReg[4]), .B(IDst[4]), .S0(ld_rec), .Y(n2630) );
  MX2X1 U2666 ( .A(IDstReg[53]), .B(IDst[53]), .S0(ld_rec), .Y(n2728) );
  MX2X1 U2667 ( .A(IDstReg[52]), .B(IDst[52]), .S0(ld_rec), .Y(n2726) );
  MX2X1 U2668 ( .A(IDstReg[51]), .B(IDst[51]), .S0(ld_rec), .Y(n2724) );
  MX2X1 U2669 ( .A(IDstReg[50]), .B(IDst[50]), .S0(ld_rec), .Y(n2722) );
  MX2X1 U2670 ( .A(IDstReg[49]), .B(IDst[49]), .S0(ld_rec), .Y(n2720) );
  OAI21X1 U2671 ( .A0(n2064), .A1(n2092), .B0(n949), .Y(DONE) );
  CLKNAND2X2 U2672 ( .A(n1243), .B(n2064), .Y(n949) );
  NOR2X1 U2673 ( .A(n2094), .B(Inst_forkAE_CONST_ENC_2_), .Y(n1243) );
  NAND4X1 U2674 ( .A(n180), .B(n179), .C(n181), .D(n2104), .Y(n2094) );
  NOR3X1 U2675 ( .A(n2065), .B(Inst_forkAE_CONST_ENC_5_), .C(
        Inst_forkAE_CONST_DEC_6_), .Y(n2104) );
  CLKINVX1 U2676 ( .A(Inst_forkAE_CONST_ENC_1_), .Y(n2065) );
  NAND4X1 U2677 ( .A(n2063), .B(n2000), .C(n185), .D(n133), .Y(n2092) );
  CLKINVX1 U2678 ( .A(Inst_forkAE_CONST_ENC_2_), .Y(n185) );
  XOR2X1 U2679 ( .A(Inst_forkAE_CONST_ENC_5_), .B(Inst_forkAE_CONST_ENC_1_), 
        .Y(n2000) );
  NOR3X1 U2680 ( .A(n1768), .B(n181), .C(n132), .Y(n2063) );
  XOR2X1 U2681 ( .A(Inst_forkAE_CONST_DEC_6_), .B(n131), .Y(n1768) );
  CLKINVX1 U2682 ( .A(n184), .Y(n2064) );
  AOI21X1 U2683 ( .A0(n957), .A1(Inst_forkAE_FSM_X_state_2_), .B0(n2087), .Y(
        n184) );
  NOR2X1 U2684 ( .A(n956), .B(Inst_forkAE_FSM_X_state_2_), .Y(n2087) );
  CLKINVX1 U2685 ( .A(Inst_forkAE_FSM_X_state_1_), .Y(n956) );
  CLKINVX1 U2686 ( .A(Inst_forkAE_FSM_X_state_0_), .Y(n957) );
endmodule

